// This is the unpowered netlist.
module sid_top (DAC_clk,
    DAC_dat_1,
    DAC_dat_2,
    DAC_le,
    bus_cyc,
    bus_we,
    clk,
    rst,
    addr,
    bus_in,
    bus_out);
 output DAC_clk;
 output DAC_dat_1;
 output DAC_dat_2;
 output DAC_le;
 input bus_cyc;
 input bus_we;
 input clk;
 input rst;
 input [5:0] addr;
 input [7:0] bus_in;
 output [7:0] bus_out;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire _06504_;
 wire _06505_;
 wire _06506_;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire _06510_;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire _06520_;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire _06527_;
 wire _06528_;
 wire _06529_;
 wire _06530_;
 wire _06531_;
 wire _06532_;
 wire _06533_;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire _06551_;
 wire _06552_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire _06557_;
 wire _06558_;
 wire _06559_;
 wire _06560_;
 wire _06561_;
 wire _06562_;
 wire _06563_;
 wire _06564_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06569_;
 wire _06570_;
 wire _06571_;
 wire _06572_;
 wire _06573_;
 wire _06574_;
 wire _06575_;
 wire _06576_;
 wire _06577_;
 wire _06578_;
 wire _06579_;
 wire _06580_;
 wire _06581_;
 wire _06582_;
 wire _06583_;
 wire _06584_;
 wire _06585_;
 wire _06586_;
 wire _06587_;
 wire _06588_;
 wire _06589_;
 wire _06590_;
 wire _06591_;
 wire _06592_;
 wire _06593_;
 wire _06594_;
 wire _06595_;
 wire _06596_;
 wire _06597_;
 wire _06598_;
 wire _06599_;
 wire _06600_;
 wire _06601_;
 wire _06602_;
 wire _06603_;
 wire _06604_;
 wire _06605_;
 wire _06606_;
 wire _06607_;
 wire _06608_;
 wire _06609_;
 wire _06610_;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire _06614_;
 wire _06615_;
 wire _06616_;
 wire _06617_;
 wire _06618_;
 wire _06619_;
 wire _06620_;
 wire _06621_;
 wire _06622_;
 wire _06623_;
 wire _06624_;
 wire _06625_;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire _06629_;
 wire _06630_;
 wire _06631_;
 wire _06632_;
 wire _06633_;
 wire _06634_;
 wire _06635_;
 wire _06636_;
 wire _06637_;
 wire _06638_;
 wire _06639_;
 wire _06640_;
 wire _06641_;
 wire _06642_;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire _06646_;
 wire _06647_;
 wire _06648_;
 wire _06649_;
 wire _06650_;
 wire _06651_;
 wire _06652_;
 wire _06653_;
 wire _06654_;
 wire _06655_;
 wire _06656_;
 wire _06657_;
 wire _06658_;
 wire _06659_;
 wire _06660_;
 wire _06661_;
 wire _06662_;
 wire _06663_;
 wire _06664_;
 wire _06665_;
 wire _06666_;
 wire _06667_;
 wire _06668_;
 wire _06669_;
 wire _06670_;
 wire _06671_;
 wire _06672_;
 wire _06673_;
 wire _06674_;
 wire _06675_;
 wire _06676_;
 wire _06677_;
 wire _06678_;
 wire _06679_;
 wire _06680_;
 wire _06681_;
 wire _06682_;
 wire _06683_;
 wire _06684_;
 wire _06685_;
 wire _06686_;
 wire _06687_;
 wire _06688_;
 wire _06689_;
 wire _06690_;
 wire _06691_;
 wire _06692_;
 wire _06693_;
 wire _06694_;
 wire _06695_;
 wire _06696_;
 wire _06697_;
 wire _06698_;
 wire _06699_;
 wire _06700_;
 wire _06701_;
 wire _06702_;
 wire _06703_;
 wire _06704_;
 wire _06705_;
 wire _06706_;
 wire _06707_;
 wire _06708_;
 wire _06709_;
 wire _06710_;
 wire _06711_;
 wire _06712_;
 wire _06713_;
 wire _06714_;
 wire _06715_;
 wire _06716_;
 wire _06717_;
 wire _06718_;
 wire _06719_;
 wire _06720_;
 wire _06721_;
 wire _06722_;
 wire _06723_;
 wire _06724_;
 wire _06725_;
 wire _06726_;
 wire _06727_;
 wire _06728_;
 wire _06729_;
 wire _06730_;
 wire _06731_;
 wire _06732_;
 wire _06733_;
 wire _06734_;
 wire _06735_;
 wire _06736_;
 wire _06737_;
 wire _06738_;
 wire _06739_;
 wire _06740_;
 wire _06741_;
 wire _06742_;
 wire _06743_;
 wire _06744_;
 wire _06745_;
 wire _06746_;
 wire _06747_;
 wire _06748_;
 wire _06749_;
 wire _06750_;
 wire _06751_;
 wire _06752_;
 wire _06753_;
 wire _06754_;
 wire _06755_;
 wire _06756_;
 wire _06757_;
 wire _06758_;
 wire _06759_;
 wire _06760_;
 wire _06761_;
 wire _06762_;
 wire _06763_;
 wire _06764_;
 wire _06765_;
 wire _06766_;
 wire _06767_;
 wire _06768_;
 wire _06769_;
 wire _06770_;
 wire _06771_;
 wire _06772_;
 wire _06773_;
 wire _06774_;
 wire _06775_;
 wire _06776_;
 wire _06777_;
 wire _06778_;
 wire _06779_;
 wire _06780_;
 wire _06781_;
 wire _06782_;
 wire _06783_;
 wire _06784_;
 wire _06785_;
 wire _06786_;
 wire _06787_;
 wire _06788_;
 wire _06789_;
 wire _06790_;
 wire _06791_;
 wire _06792_;
 wire _06793_;
 wire _06794_;
 wire _06795_;
 wire _06796_;
 wire _06797_;
 wire _06798_;
 wire _06799_;
 wire _06800_;
 wire _06801_;
 wire _06802_;
 wire _06803_;
 wire _06804_;
 wire _06805_;
 wire _06806_;
 wire _06807_;
 wire _06808_;
 wire _06809_;
 wire _06810_;
 wire _06811_;
 wire _06812_;
 wire _06813_;
 wire _06814_;
 wire _06815_;
 wire _06816_;
 wire _06817_;
 wire _06818_;
 wire _06819_;
 wire _06820_;
 wire _06821_;
 wire _06822_;
 wire _06823_;
 wire _06824_;
 wire _06825_;
 wire _06826_;
 wire _06827_;
 wire _06828_;
 wire _06829_;
 wire _06830_;
 wire _06831_;
 wire _06832_;
 wire _06833_;
 wire _06834_;
 wire _06835_;
 wire _06836_;
 wire _06837_;
 wire _06838_;
 wire _06839_;
 wire _06840_;
 wire _06841_;
 wire _06842_;
 wire _06843_;
 wire _06844_;
 wire _06845_;
 wire _06846_;
 wire _06847_;
 wire _06848_;
 wire _06849_;
 wire _06850_;
 wire _06851_;
 wire _06852_;
 wire _06853_;
 wire _06854_;
 wire _06855_;
 wire _06856_;
 wire _06857_;
 wire _06858_;
 wire _06859_;
 wire _06860_;
 wire _06861_;
 wire _06862_;
 wire _06863_;
 wire _06864_;
 wire _06865_;
 wire _06866_;
 wire _06867_;
 wire _06868_;
 wire _06869_;
 wire _06870_;
 wire _06871_;
 wire _06872_;
 wire _06873_;
 wire _06874_;
 wire _06875_;
 wire _06876_;
 wire _06877_;
 wire _06878_;
 wire _06879_;
 wire _06880_;
 wire _06881_;
 wire _06882_;
 wire _06883_;
 wire _06884_;
 wire _06885_;
 wire _06886_;
 wire _06887_;
 wire _06888_;
 wire _06889_;
 wire _06890_;
 wire _06891_;
 wire _06892_;
 wire _06893_;
 wire _06894_;
 wire _06895_;
 wire _06896_;
 wire _06897_;
 wire _06898_;
 wire _06899_;
 wire _06900_;
 wire _06901_;
 wire _06902_;
 wire _06903_;
 wire _06904_;
 wire _06905_;
 wire _06906_;
 wire _06907_;
 wire _06908_;
 wire _06909_;
 wire _06910_;
 wire _06911_;
 wire _06912_;
 wire _06913_;
 wire _06914_;
 wire _06915_;
 wire _06916_;
 wire _06917_;
 wire _06918_;
 wire _06919_;
 wire _06920_;
 wire _06921_;
 wire _06922_;
 wire _06923_;
 wire _06924_;
 wire _06925_;
 wire _06926_;
 wire _06927_;
 wire _06928_;
 wire _06929_;
 wire _06930_;
 wire _06931_;
 wire _06932_;
 wire _06933_;
 wire _06934_;
 wire _06935_;
 wire _06936_;
 wire _06937_;
 wire _06938_;
 wire _06939_;
 wire _06940_;
 wire _06941_;
 wire _06942_;
 wire _06943_;
 wire _06944_;
 wire _06945_;
 wire _06946_;
 wire _06947_;
 wire _06948_;
 wire _06949_;
 wire _06950_;
 wire _06951_;
 wire _06952_;
 wire _06953_;
 wire _06954_;
 wire _06955_;
 wire _06956_;
 wire _06957_;
 wire _06958_;
 wire _06959_;
 wire _06960_;
 wire _06961_;
 wire _06962_;
 wire _06963_;
 wire _06964_;
 wire _06965_;
 wire _06966_;
 wire _06967_;
 wire _06968_;
 wire _06969_;
 wire _06970_;
 wire _06971_;
 wire _06972_;
 wire _06973_;
 wire _06974_;
 wire _06975_;
 wire _06976_;
 wire _06977_;
 wire _06978_;
 wire _06979_;
 wire _06980_;
 wire _06981_;
 wire _06982_;
 wire _06983_;
 wire _06984_;
 wire _06985_;
 wire _06986_;
 wire _06987_;
 wire _06988_;
 wire _06989_;
 wire _06990_;
 wire _06991_;
 wire _06992_;
 wire _06993_;
 wire _06994_;
 wire _06995_;
 wire _06996_;
 wire _06997_;
 wire _06998_;
 wire _06999_;
 wire _07000_;
 wire _07001_;
 wire _07002_;
 wire _07003_;
 wire _07004_;
 wire _07005_;
 wire _07006_;
 wire _07007_;
 wire _07008_;
 wire _07009_;
 wire _07010_;
 wire _07011_;
 wire _07012_;
 wire _07013_;
 wire _07014_;
 wire _07015_;
 wire _07016_;
 wire _07017_;
 wire _07018_;
 wire _07019_;
 wire _07020_;
 wire _07021_;
 wire _07022_;
 wire _07023_;
 wire _07024_;
 wire _07025_;
 wire _07026_;
 wire _07027_;
 wire _07028_;
 wire _07029_;
 wire _07030_;
 wire _07031_;
 wire _07032_;
 wire _07033_;
 wire _07034_;
 wire _07035_;
 wire _07036_;
 wire _07037_;
 wire _07038_;
 wire _07039_;
 wire _07040_;
 wire _07041_;
 wire _07042_;
 wire _07043_;
 wire _07044_;
 wire _07045_;
 wire _07046_;
 wire _07047_;
 wire _07048_;
 wire _07049_;
 wire _07050_;
 wire _07051_;
 wire _07052_;
 wire _07053_;
 wire _07054_;
 wire _07055_;
 wire _07056_;
 wire _07057_;
 wire _07058_;
 wire _07059_;
 wire _07060_;
 wire _07061_;
 wire _07062_;
 wire _07063_;
 wire _07064_;
 wire _07065_;
 wire _07066_;
 wire _07067_;
 wire _07068_;
 wire _07069_;
 wire _07070_;
 wire _07071_;
 wire _07072_;
 wire _07073_;
 wire _07074_;
 wire _07075_;
 wire _07076_;
 wire _07077_;
 wire _07078_;
 wire _07079_;
 wire _07080_;
 wire _07081_;
 wire _07082_;
 wire _07083_;
 wire _07084_;
 wire _07085_;
 wire _07086_;
 wire _07087_;
 wire _07088_;
 wire _07089_;
 wire _07090_;
 wire _07091_;
 wire _07092_;
 wire _07093_;
 wire _07094_;
 wire _07095_;
 wire _07096_;
 wire _07097_;
 wire _07098_;
 wire _07099_;
 wire _07100_;
 wire _07101_;
 wire _07102_;
 wire _07103_;
 wire _07104_;
 wire _07105_;
 wire _07106_;
 wire _07107_;
 wire _07108_;
 wire _07109_;
 wire _07110_;
 wire _07111_;
 wire _07112_;
 wire _07113_;
 wire _07114_;
 wire _07115_;
 wire _07116_;
 wire _07117_;
 wire _07118_;
 wire _07119_;
 wire _07120_;
 wire _07121_;
 wire _07122_;
 wire _07123_;
 wire _07124_;
 wire _07125_;
 wire _07126_;
 wire _07127_;
 wire _07128_;
 wire _07129_;
 wire _07130_;
 wire _07131_;
 wire _07132_;
 wire _07133_;
 wire _07134_;
 wire _07135_;
 wire _07136_;
 wire _07137_;
 wire _07138_;
 wire _07139_;
 wire _07140_;
 wire _07141_;
 wire _07142_;
 wire _07143_;
 wire _07144_;
 wire _07145_;
 wire _07146_;
 wire _07147_;
 wire _07148_;
 wire _07149_;
 wire _07150_;
 wire _07151_;
 wire _07152_;
 wire _07153_;
 wire _07154_;
 wire _07155_;
 wire _07156_;
 wire _07157_;
 wire _07158_;
 wire _07159_;
 wire _07160_;
 wire _07161_;
 wire _07162_;
 wire _07163_;
 wire _07164_;
 wire _07165_;
 wire _07166_;
 wire _07167_;
 wire _07168_;
 wire _07169_;
 wire _07170_;
 wire _07171_;
 wire _07172_;
 wire _07173_;
 wire _07174_;
 wire _07175_;
 wire _07176_;
 wire _07177_;
 wire _07178_;
 wire _07179_;
 wire _07180_;
 wire _07181_;
 wire _07182_;
 wire _07183_;
 wire _07184_;
 wire _07185_;
 wire _07186_;
 wire _07187_;
 wire _07188_;
 wire _07189_;
 wire _07190_;
 wire _07191_;
 wire _07192_;
 wire _07193_;
 wire _07194_;
 wire _07195_;
 wire _07196_;
 wire _07197_;
 wire _07198_;
 wire _07199_;
 wire _07200_;
 wire _07201_;
 wire _07202_;
 wire _07203_;
 wire _07204_;
 wire _07205_;
 wire _07206_;
 wire _07207_;
 wire _07208_;
 wire _07209_;
 wire _07210_;
 wire _07211_;
 wire _07212_;
 wire _07213_;
 wire _07214_;
 wire _07215_;
 wire _07216_;
 wire _07217_;
 wire _07218_;
 wire _07219_;
 wire _07220_;
 wire _07221_;
 wire _07222_;
 wire _07223_;
 wire _07224_;
 wire _07225_;
 wire _07226_;
 wire _07227_;
 wire _07228_;
 wire _07229_;
 wire _07230_;
 wire _07231_;
 wire _07232_;
 wire _07233_;
 wire _07234_;
 wire _07235_;
 wire _07236_;
 wire _07237_;
 wire _07238_;
 wire _07239_;
 wire _07240_;
 wire _07241_;
 wire _07242_;
 wire _07243_;
 wire _07244_;
 wire _07245_;
 wire _07246_;
 wire _07247_;
 wire _07248_;
 wire _07249_;
 wire _07250_;
 wire _07251_;
 wire _07252_;
 wire _07253_;
 wire _07254_;
 wire _07255_;
 wire _07256_;
 wire _07257_;
 wire _07258_;
 wire _07259_;
 wire _07260_;
 wire _07261_;
 wire _07262_;
 wire _07263_;
 wire _07264_;
 wire _07265_;
 wire _07266_;
 wire _07267_;
 wire _07268_;
 wire _07269_;
 wire _07270_;
 wire _07271_;
 wire _07272_;
 wire _07273_;
 wire _07274_;
 wire _07275_;
 wire _07276_;
 wire _07277_;
 wire _07278_;
 wire _07279_;
 wire _07280_;
 wire _07281_;
 wire _07282_;
 wire _07283_;
 wire _07284_;
 wire _07285_;
 wire _07286_;
 wire _07287_;
 wire _07288_;
 wire _07289_;
 wire _07290_;
 wire _07291_;
 wire _07292_;
 wire _07293_;
 wire _07294_;
 wire _07295_;
 wire _07296_;
 wire _07297_;
 wire _07298_;
 wire _07299_;
 wire _07300_;
 wire _07301_;
 wire _07302_;
 wire _07303_;
 wire _07304_;
 wire _07305_;
 wire _07306_;
 wire _07307_;
 wire _07308_;
 wire _07309_;
 wire _07310_;
 wire _07311_;
 wire _07312_;
 wire _07313_;
 wire _07314_;
 wire _07315_;
 wire _07316_;
 wire _07317_;
 wire _07318_;
 wire _07319_;
 wire _07320_;
 wire _07321_;
 wire _07322_;
 wire _07323_;
 wire _07324_;
 wire _07325_;
 wire _07326_;
 wire _07327_;
 wire _07328_;
 wire _07329_;
 wire _07330_;
 wire _07331_;
 wire _07332_;
 wire _07333_;
 wire _07334_;
 wire _07335_;
 wire _07336_;
 wire _07337_;
 wire _07338_;
 wire _07339_;
 wire _07340_;
 wire _07341_;
 wire _07342_;
 wire _07343_;
 wire _07344_;
 wire _07345_;
 wire _07346_;
 wire _07347_;
 wire _07348_;
 wire _07349_;
 wire _07350_;
 wire _07351_;
 wire _07352_;
 wire _07353_;
 wire _07354_;
 wire _07355_;
 wire _07356_;
 wire _07357_;
 wire _07358_;
 wire _07359_;
 wire _07360_;
 wire _07361_;
 wire _07362_;
 wire _07363_;
 wire _07364_;
 wire _07365_;
 wire _07366_;
 wire _07367_;
 wire _07368_;
 wire _07369_;
 wire _07370_;
 wire _07371_;
 wire _07372_;
 wire _07373_;
 wire _07374_;
 wire _07375_;
 wire _07376_;
 wire _07377_;
 wire _07378_;
 wire _07379_;
 wire _07380_;
 wire _07381_;
 wire _07382_;
 wire _07383_;
 wire _07384_;
 wire _07385_;
 wire _07386_;
 wire _07387_;
 wire _07388_;
 wire _07389_;
 wire _07390_;
 wire _07391_;
 wire _07392_;
 wire _07393_;
 wire _07394_;
 wire _07395_;
 wire _07396_;
 wire _07397_;
 wire _07398_;
 wire _07399_;
 wire _07400_;
 wire _07401_;
 wire _07402_;
 wire _07403_;
 wire _07404_;
 wire _07405_;
 wire _07406_;
 wire _07407_;
 wire _07408_;
 wire _07409_;
 wire _07410_;
 wire _07411_;
 wire _07412_;
 wire _07413_;
 wire _07414_;
 wire _07415_;
 wire _07416_;
 wire _07417_;
 wire _07418_;
 wire _07419_;
 wire _07420_;
 wire _07421_;
 wire _07422_;
 wire _07423_;
 wire _07424_;
 wire _07425_;
 wire _07426_;
 wire _07427_;
 wire _07428_;
 wire _07429_;
 wire _07430_;
 wire _07431_;
 wire _07432_;
 wire _07433_;
 wire _07434_;
 wire _07435_;
 wire _07436_;
 wire _07437_;
 wire _07438_;
 wire _07439_;
 wire _07440_;
 wire _07441_;
 wire _07442_;
 wire _07443_;
 wire _07444_;
 wire _07445_;
 wire _07446_;
 wire _07447_;
 wire _07448_;
 wire _07449_;
 wire _07450_;
 wire _07451_;
 wire _07452_;
 wire _07453_;
 wire _07454_;
 wire _07455_;
 wire _07456_;
 wire _07457_;
 wire _07458_;
 wire _07459_;
 wire _07460_;
 wire _07461_;
 wire _07462_;
 wire _07463_;
 wire _07464_;
 wire _07465_;
 wire _07466_;
 wire _07467_;
 wire _07468_;
 wire _07469_;
 wire _07470_;
 wire _07471_;
 wire _07472_;
 wire _07473_;
 wire _07474_;
 wire _07475_;
 wire _07476_;
 wire _07477_;
 wire _07478_;
 wire _07479_;
 wire _07480_;
 wire _07481_;
 wire _07482_;
 wire _07483_;
 wire _07484_;
 wire _07485_;
 wire _07486_;
 wire _07487_;
 wire _07488_;
 wire _07489_;
 wire _07490_;
 wire _07491_;
 wire _07492_;
 wire _07493_;
 wire _07494_;
 wire _07495_;
 wire _07496_;
 wire _07497_;
 wire _07498_;
 wire _07499_;
 wire _07500_;
 wire _07501_;
 wire _07502_;
 wire _07503_;
 wire _07504_;
 wire _07505_;
 wire _07506_;
 wire _07507_;
 wire _07508_;
 wire _07509_;
 wire _07510_;
 wire _07511_;
 wire _07512_;
 wire _07513_;
 wire _07514_;
 wire _07515_;
 wire _07516_;
 wire _07517_;
 wire _07518_;
 wire _07519_;
 wire _07520_;
 wire _07521_;
 wire _07522_;
 wire _07523_;
 wire _07524_;
 wire _07525_;
 wire _07526_;
 wire _07527_;
 wire _07528_;
 wire _07529_;
 wire _07530_;
 wire _07531_;
 wire _07532_;
 wire _07533_;
 wire _07534_;
 wire _07535_;
 wire _07536_;
 wire _07537_;
 wire _07538_;
 wire _07539_;
 wire _07540_;
 wire _07541_;
 wire _07542_;
 wire _07543_;
 wire _07544_;
 wire _07545_;
 wire _07546_;
 wire _07547_;
 wire _07548_;
 wire _07549_;
 wire _07550_;
 wire _07551_;
 wire _07552_;
 wire _07553_;
 wire _07554_;
 wire _07555_;
 wire _07556_;
 wire _07557_;
 wire _07558_;
 wire _07559_;
 wire _07560_;
 wire _07561_;
 wire _07562_;
 wire _07563_;
 wire _07564_;
 wire _07565_;
 wire _07566_;
 wire _07567_;
 wire _07568_;
 wire _07569_;
 wire _07570_;
 wire _07571_;
 wire _07572_;
 wire _07573_;
 wire _07574_;
 wire _07575_;
 wire _07576_;
 wire _07577_;
 wire _07578_;
 wire _07579_;
 wire _07580_;
 wire _07581_;
 wire _07582_;
 wire _07583_;
 wire _07584_;
 wire _07585_;
 wire _07586_;
 wire _07587_;
 wire _07588_;
 wire _07589_;
 wire _07590_;
 wire _07591_;
 wire _07592_;
 wire _07593_;
 wire _07594_;
 wire _07595_;
 wire _07596_;
 wire _07597_;
 wire _07598_;
 wire _07599_;
 wire _07600_;
 wire _07601_;
 wire _07602_;
 wire _07603_;
 wire _07604_;
 wire _07605_;
 wire _07606_;
 wire _07607_;
 wire _07608_;
 wire _07609_;
 wire _07610_;
 wire _07611_;
 wire _07612_;
 wire _07613_;
 wire _07614_;
 wire _07615_;
 wire _07616_;
 wire _07617_;
 wire _07618_;
 wire _07619_;
 wire _07620_;
 wire _07621_;
 wire _07622_;
 wire _07623_;
 wire _07624_;
 wire _07625_;
 wire _07626_;
 wire _07627_;
 wire _07628_;
 wire _07629_;
 wire _07630_;
 wire _07631_;
 wire _07632_;
 wire _07633_;
 wire _07634_;
 wire _07635_;
 wire _07636_;
 wire _07637_;
 wire _07638_;
 wire _07639_;
 wire _07640_;
 wire _07641_;
 wire _07642_;
 wire _07643_;
 wire _07644_;
 wire _07645_;
 wire _07646_;
 wire _07647_;
 wire _07648_;
 wire _07649_;
 wire _07650_;
 wire _07651_;
 wire _07652_;
 wire _07653_;
 wire _07654_;
 wire _07655_;
 wire _07656_;
 wire _07657_;
 wire _07658_;
 wire _07659_;
 wire _07660_;
 wire _07661_;
 wire _07662_;
 wire _07663_;
 wire _07664_;
 wire _07665_;
 wire _07666_;
 wire _07667_;
 wire _07668_;
 wire _07669_;
 wire _07670_;
 wire _07671_;
 wire _07672_;
 wire _07673_;
 wire _07674_;
 wire _07675_;
 wire _07676_;
 wire _07677_;
 wire _07678_;
 wire _07679_;
 wire _07680_;
 wire _07681_;
 wire _07682_;
 wire _07683_;
 wire _07684_;
 wire _07685_;
 wire _07686_;
 wire _07687_;
 wire _07688_;
 wire _07689_;
 wire _07690_;
 wire _07691_;
 wire _07692_;
 wire _07693_;
 wire _07694_;
 wire _07695_;
 wire _07696_;
 wire _07697_;
 wire _07698_;
 wire _07699_;
 wire _07700_;
 wire _07701_;
 wire _07702_;
 wire _07703_;
 wire _07704_;
 wire _07705_;
 wire _07706_;
 wire _07707_;
 wire _07708_;
 wire _07709_;
 wire _07710_;
 wire _07711_;
 wire _07712_;
 wire _07713_;
 wire _07714_;
 wire _07715_;
 wire _07716_;
 wire _07717_;
 wire _07718_;
 wire _07719_;
 wire _07720_;
 wire _07721_;
 wire _07722_;
 wire _07723_;
 wire _07724_;
 wire _07725_;
 wire _07726_;
 wire _07727_;
 wire _07728_;
 wire _07729_;
 wire _07730_;
 wire _07731_;
 wire _07732_;
 wire _07733_;
 wire _07734_;
 wire _07735_;
 wire _07736_;
 wire _07737_;
 wire _07738_;
 wire _07739_;
 wire _07740_;
 wire _07741_;
 wire _07742_;
 wire _07743_;
 wire _07744_;
 wire _07745_;
 wire _07746_;
 wire _07747_;
 wire _07748_;
 wire _07749_;
 wire _07750_;
 wire _07751_;
 wire _07752_;
 wire _07753_;
 wire _07754_;
 wire _07755_;
 wire _07756_;
 wire _07757_;
 wire _07758_;
 wire _07759_;
 wire _07760_;
 wire _07761_;
 wire _07762_;
 wire _07763_;
 wire _07764_;
 wire _07765_;
 wire _07766_;
 wire _07767_;
 wire _07768_;
 wire _07769_;
 wire _07770_;
 wire _07771_;
 wire _07772_;
 wire _07773_;
 wire _07774_;
 wire _07775_;
 wire _07776_;
 wire _07777_;
 wire _07778_;
 wire _07779_;
 wire _07780_;
 wire _07781_;
 wire _07782_;
 wire _07783_;
 wire _07784_;
 wire _07785_;
 wire _07786_;
 wire _07787_;
 wire _07788_;
 wire _07789_;
 wire _07790_;
 wire _07791_;
 wire _07792_;
 wire _07793_;
 wire _07794_;
 wire _07795_;
 wire _07796_;
 wire _07797_;
 wire _07798_;
 wire _07799_;
 wire _07800_;
 wire _07801_;
 wire _07802_;
 wire _07803_;
 wire _07804_;
 wire _07805_;
 wire _07806_;
 wire _07807_;
 wire _07808_;
 wire _07809_;
 wire _07810_;
 wire _07811_;
 wire _07812_;
 wire _07813_;
 wire _07814_;
 wire _07815_;
 wire _07816_;
 wire _07817_;
 wire _07818_;
 wire _07819_;
 wire _07820_;
 wire _07821_;
 wire _07822_;
 wire _07823_;
 wire _07824_;
 wire _07825_;
 wire _07826_;
 wire _07827_;
 wire _07828_;
 wire _07829_;
 wire _07830_;
 wire _07831_;
 wire _07832_;
 wire _07833_;
 wire _07834_;
 wire _07835_;
 wire _07836_;
 wire _07837_;
 wire _07838_;
 wire _07839_;
 wire _07840_;
 wire _07841_;
 wire _07842_;
 wire _07843_;
 wire _07844_;
 wire _07845_;
 wire _07846_;
 wire _07847_;
 wire _07848_;
 wire _07849_;
 wire _07850_;
 wire _07851_;
 wire _07852_;
 wire _07853_;
 wire _07854_;
 wire _07855_;
 wire _07856_;
 wire _07857_;
 wire _07858_;
 wire _07859_;
 wire _07860_;
 wire _07861_;
 wire _07862_;
 wire _07863_;
 wire _07864_;
 wire _07865_;
 wire _07866_;
 wire _07867_;
 wire _07868_;
 wire _07869_;
 wire _07870_;
 wire _07871_;
 wire _07872_;
 wire _07873_;
 wire _07874_;
 wire _07875_;
 wire _07876_;
 wire _07877_;
 wire _07878_;
 wire _07879_;
 wire _07880_;
 wire _07881_;
 wire _07882_;
 wire _07883_;
 wire _07884_;
 wire _07885_;
 wire _07886_;
 wire _07887_;
 wire _07888_;
 wire _07889_;
 wire _07890_;
 wire _07891_;
 wire _07892_;
 wire _07893_;
 wire _07894_;
 wire _07895_;
 wire _07896_;
 wire _07897_;
 wire _07898_;
 wire _07899_;
 wire _07900_;
 wire _07901_;
 wire _07902_;
 wire _07903_;
 wire _07904_;
 wire _07905_;
 wire _07906_;
 wire _07907_;
 wire _07908_;
 wire _07909_;
 wire _07910_;
 wire _07911_;
 wire _07912_;
 wire _07913_;
 wire _07914_;
 wire _07915_;
 wire _07916_;
 wire _07917_;
 wire _07918_;
 wire _07919_;
 wire _07920_;
 wire _07921_;
 wire _07922_;
 wire _07923_;
 wire _07924_;
 wire _07925_;
 wire _07926_;
 wire _07927_;
 wire _07928_;
 wire _07929_;
 wire _07930_;
 wire _07931_;
 wire _07932_;
 wire _07933_;
 wire _07934_;
 wire _07935_;
 wire _07936_;
 wire _07937_;
 wire _07938_;
 wire _07939_;
 wire _07940_;
 wire _07941_;
 wire _07942_;
 wire _07943_;
 wire _07944_;
 wire _07945_;
 wire _07946_;
 wire _07947_;
 wire _07948_;
 wire _07949_;
 wire _07950_;
 wire _07951_;
 wire _07952_;
 wire _07953_;
 wire _07954_;
 wire _07955_;
 wire _07956_;
 wire _07957_;
 wire _07958_;
 wire _07959_;
 wire _07960_;
 wire _07961_;
 wire _07962_;
 wire _07963_;
 wire _07964_;
 wire _07965_;
 wire _07966_;
 wire _07967_;
 wire _07968_;
 wire _07969_;
 wire _07970_;
 wire _07971_;
 wire _07972_;
 wire _07973_;
 wire _07974_;
 wire _07975_;
 wire _07976_;
 wire _07977_;
 wire _07978_;
 wire _07979_;
 wire _07980_;
 wire _07981_;
 wire _07982_;
 wire _07983_;
 wire _07984_;
 wire _07985_;
 wire _07986_;
 wire _07987_;
 wire _07988_;
 wire _07989_;
 wire _07990_;
 wire _07991_;
 wire _07992_;
 wire _07993_;
 wire _07994_;
 wire _07995_;
 wire _07996_;
 wire _07997_;
 wire _07998_;
 wire _07999_;
 wire _08000_;
 wire _08001_;
 wire _08002_;
 wire _08003_;
 wire _08004_;
 wire _08005_;
 wire _08006_;
 wire _08007_;
 wire _08008_;
 wire _08009_;
 wire _08010_;
 wire _08011_;
 wire _08012_;
 wire _08013_;
 wire _08014_;
 wire _08015_;
 wire _08016_;
 wire _08017_;
 wire _08018_;
 wire _08019_;
 wire _08020_;
 wire _08021_;
 wire _08022_;
 wire _08023_;
 wire _08024_;
 wire _08025_;
 wire _08026_;
 wire _08027_;
 wire _08028_;
 wire _08029_;
 wire _08030_;
 wire _08031_;
 wire _08032_;
 wire _08033_;
 wire _08034_;
 wire _08035_;
 wire _08036_;
 wire _08037_;
 wire _08038_;
 wire _08039_;
 wire _08040_;
 wire _08041_;
 wire _08042_;
 wire _08043_;
 wire _08044_;
 wire _08045_;
 wire _08046_;
 wire _08047_;
 wire _08048_;
 wire _08049_;
 wire _08050_;
 wire _08051_;
 wire _08052_;
 wire _08053_;
 wire _08054_;
 wire _08055_;
 wire _08056_;
 wire _08057_;
 wire _08058_;
 wire _08059_;
 wire _08060_;
 wire _08061_;
 wire _08062_;
 wire _08063_;
 wire _08064_;
 wire _08065_;
 wire _08066_;
 wire _08067_;
 wire _08068_;
 wire _08069_;
 wire _08070_;
 wire _08071_;
 wire _08072_;
 wire _08073_;
 wire _08074_;
 wire _08075_;
 wire _08076_;
 wire _08077_;
 wire _08078_;
 wire _08079_;
 wire _08080_;
 wire _08081_;
 wire _08082_;
 wire _08083_;
 wire _08084_;
 wire _08085_;
 wire _08086_;
 wire _08087_;
 wire _08088_;
 wire _08089_;
 wire _08090_;
 wire _08091_;
 wire _08092_;
 wire _08093_;
 wire _08094_;
 wire _08095_;
 wire _08096_;
 wire _08097_;
 wire _08098_;
 wire _08099_;
 wire _08100_;
 wire _08101_;
 wire _08102_;
 wire _08103_;
 wire _08104_;
 wire _08105_;
 wire _08106_;
 wire _08107_;
 wire _08108_;
 wire _08109_;
 wire _08110_;
 wire _08111_;
 wire _08112_;
 wire _08113_;
 wire _08114_;
 wire _08115_;
 wire _08116_;
 wire _08117_;
 wire _08118_;
 wire _08119_;
 wire _08120_;
 wire _08121_;
 wire _08122_;
 wire _08123_;
 wire _08124_;
 wire _08125_;
 wire _08126_;
 wire _08127_;
 wire _08128_;
 wire _08129_;
 wire _08130_;
 wire _08131_;
 wire _08132_;
 wire _08133_;
 wire _08134_;
 wire _08135_;
 wire _08136_;
 wire _08137_;
 wire _08138_;
 wire _08139_;
 wire _08140_;
 wire _08141_;
 wire _08142_;
 wire _08143_;
 wire _08144_;
 wire _08145_;
 wire _08146_;
 wire _08147_;
 wire _08148_;
 wire _08149_;
 wire _08150_;
 wire _08151_;
 wire _08152_;
 wire _08153_;
 wire _08154_;
 wire _08155_;
 wire _08156_;
 wire _08157_;
 wire _08158_;
 wire _08159_;
 wire _08160_;
 wire _08161_;
 wire _08162_;
 wire _08163_;
 wire _08164_;
 wire _08165_;
 wire _08166_;
 wire _08167_;
 wire _08168_;
 wire _08169_;
 wire _08170_;
 wire _08171_;
 wire _08172_;
 wire _08173_;
 wire _08174_;
 wire _08175_;
 wire _08176_;
 wire _08177_;
 wire _08178_;
 wire _08179_;
 wire _08180_;
 wire _08181_;
 wire _08182_;
 wire _08183_;
 wire _08184_;
 wire _08185_;
 wire _08186_;
 wire _08187_;
 wire _08188_;
 wire _08189_;
 wire _08190_;
 wire _08191_;
 wire _08192_;
 wire _08193_;
 wire _08194_;
 wire _08195_;
 wire _08196_;
 wire _08197_;
 wire _08198_;
 wire _08199_;
 wire _08200_;
 wire _08201_;
 wire _08202_;
 wire _08203_;
 wire _08204_;
 wire _08205_;
 wire _08206_;
 wire _08207_;
 wire _08208_;
 wire _08209_;
 wire _08210_;
 wire _08211_;
 wire _08212_;
 wire _08213_;
 wire _08214_;
 wire _08215_;
 wire _08216_;
 wire _08217_;
 wire _08218_;
 wire _08219_;
 wire _08220_;
 wire _08221_;
 wire _08222_;
 wire _08223_;
 wire _08224_;
 wire _08225_;
 wire _08226_;
 wire _08227_;
 wire _08228_;
 wire _08229_;
 wire _08230_;
 wire _08231_;
 wire _08232_;
 wire _08233_;
 wire _08234_;
 wire _08235_;
 wire _08236_;
 wire _08237_;
 wire _08238_;
 wire _08239_;
 wire _08240_;
 wire _08241_;
 wire _08242_;
 wire _08243_;
 wire _08244_;
 wire _08245_;
 wire _08246_;
 wire _08247_;
 wire _08248_;
 wire _08249_;
 wire _08250_;
 wire _08251_;
 wire _08252_;
 wire _08253_;
 wire _08254_;
 wire _08255_;
 wire _08256_;
 wire _08257_;
 wire _08258_;
 wire _08259_;
 wire _08260_;
 wire _08261_;
 wire _08262_;
 wire _08263_;
 wire _08264_;
 wire _08265_;
 wire _08266_;
 wire _08267_;
 wire _08268_;
 wire _08269_;
 wire _08270_;
 wire _08271_;
 wire _08272_;
 wire _08273_;
 wire _08274_;
 wire _08275_;
 wire _08276_;
 wire _08277_;
 wire _08278_;
 wire _08279_;
 wire _08280_;
 wire _08281_;
 wire _08282_;
 wire _08283_;
 wire _08284_;
 wire _08285_;
 wire _08286_;
 wire _08287_;
 wire _08288_;
 wire _08289_;
 wire _08290_;
 wire _08291_;
 wire _08292_;
 wire _08293_;
 wire _08294_;
 wire _08295_;
 wire _08296_;
 wire _08297_;
 wire _08298_;
 wire _08299_;
 wire _08300_;
 wire _08301_;
 wire _08302_;
 wire _08303_;
 wire _08304_;
 wire _08305_;
 wire _08306_;
 wire _08307_;
 wire _08308_;
 wire _08309_;
 wire _08310_;
 wire _08311_;
 wire _08312_;
 wire _08313_;
 wire _08314_;
 wire _08315_;
 wire _08316_;
 wire _08317_;
 wire _08318_;
 wire _08319_;
 wire _08320_;
 wire _08321_;
 wire _08322_;
 wire _08323_;
 wire _08324_;
 wire _08325_;
 wire _08326_;
 wire _08327_;
 wire _08328_;
 wire _08329_;
 wire _08330_;
 wire _08331_;
 wire _08332_;
 wire _08333_;
 wire _08334_;
 wire _08335_;
 wire _08336_;
 wire _08337_;
 wire _08338_;
 wire _08339_;
 wire _08340_;
 wire _08341_;
 wire _08342_;
 wire _08343_;
 wire _08344_;
 wire _08345_;
 wire _08346_;
 wire _08347_;
 wire _08348_;
 wire _08349_;
 wire _08350_;
 wire _08351_;
 wire _08352_;
 wire _08353_;
 wire _08354_;
 wire _08355_;
 wire _08356_;
 wire _08357_;
 wire _08358_;
 wire _08359_;
 wire _08360_;
 wire _08361_;
 wire _08362_;
 wire _08363_;
 wire _08364_;
 wire _08365_;
 wire _08366_;
 wire _08367_;
 wire _08368_;
 wire _08369_;
 wire _08370_;
 wire _08371_;
 wire _08372_;
 wire _08373_;
 wire _08374_;
 wire _08375_;
 wire _08376_;
 wire _08377_;
 wire _08378_;
 wire _08379_;
 wire _08380_;
 wire _08381_;
 wire _08382_;
 wire _08383_;
 wire _08384_;
 wire _08385_;
 wire _08386_;
 wire _08387_;
 wire _08388_;
 wire _08389_;
 wire _08390_;
 wire _08391_;
 wire _08392_;
 wire _08393_;
 wire _08394_;
 wire _08395_;
 wire _08396_;
 wire _08397_;
 wire _08398_;
 wire _08399_;
 wire _08400_;
 wire _08401_;
 wire _08402_;
 wire _08403_;
 wire _08404_;
 wire _08405_;
 wire _08406_;
 wire _08407_;
 wire _08408_;
 wire _08409_;
 wire _08410_;
 wire _08411_;
 wire _08412_;
 wire _08413_;
 wire _08414_;
 wire _08415_;
 wire _08416_;
 wire _08417_;
 wire _08418_;
 wire _08419_;
 wire _08420_;
 wire _08421_;
 wire _08422_;
 wire _08423_;
 wire _08424_;
 wire _08425_;
 wire _08426_;
 wire _08427_;
 wire _08428_;
 wire _08429_;
 wire _08430_;
 wire _08431_;
 wire _08432_;
 wire _08433_;
 wire _08434_;
 wire _08435_;
 wire _08436_;
 wire _08437_;
 wire _08438_;
 wire _08439_;
 wire _08440_;
 wire _08441_;
 wire _08442_;
 wire _08443_;
 wire _08444_;
 wire _08445_;
 wire _08446_;
 wire _08447_;
 wire _08448_;
 wire _08449_;
 wire _08450_;
 wire _08451_;
 wire _08452_;
 wire _08453_;
 wire _08454_;
 wire _08455_;
 wire _08456_;
 wire _08457_;
 wire _08458_;
 wire _08459_;
 wire _08460_;
 wire _08461_;
 wire _08462_;
 wire _08463_;
 wire _08464_;
 wire _08465_;
 wire _08466_;
 wire \channels.accum[0][0] ;
 wire \channels.accum[0][10] ;
 wire \channels.accum[0][11] ;
 wire \channels.accum[0][12] ;
 wire \channels.accum[0][13] ;
 wire \channels.accum[0][14] ;
 wire \channels.accum[0][15] ;
 wire \channels.accum[0][16] ;
 wire \channels.accum[0][17] ;
 wire \channels.accum[0][18] ;
 wire \channels.accum[0][19] ;
 wire \channels.accum[0][1] ;
 wire \channels.accum[0][20] ;
 wire \channels.accum[0][21] ;
 wire \channels.accum[0][22] ;
 wire \channels.accum[0][23] ;
 wire \channels.accum[0][2] ;
 wire \channels.accum[0][3] ;
 wire \channels.accum[0][4] ;
 wire \channels.accum[0][5] ;
 wire \channels.accum[0][6] ;
 wire \channels.accum[0][7] ;
 wire \channels.accum[0][8] ;
 wire \channels.accum[0][9] ;
 wire \channels.accum[1][0] ;
 wire \channels.accum[1][10] ;
 wire \channels.accum[1][11] ;
 wire \channels.accum[1][12] ;
 wire \channels.accum[1][13] ;
 wire \channels.accum[1][14] ;
 wire \channels.accum[1][15] ;
 wire \channels.accum[1][16] ;
 wire \channels.accum[1][17] ;
 wire \channels.accum[1][18] ;
 wire \channels.accum[1][19] ;
 wire \channels.accum[1][1] ;
 wire \channels.accum[1][20] ;
 wire \channels.accum[1][21] ;
 wire \channels.accum[1][22] ;
 wire \channels.accum[1][23] ;
 wire \channels.accum[1][2] ;
 wire \channels.accum[1][3] ;
 wire \channels.accum[1][4] ;
 wire \channels.accum[1][5] ;
 wire \channels.accum[1][6] ;
 wire \channels.accum[1][7] ;
 wire \channels.accum[1][8] ;
 wire \channels.accum[1][9] ;
 wire \channels.accum[2][0] ;
 wire \channels.accum[2][10] ;
 wire \channels.accum[2][11] ;
 wire \channels.accum[2][12] ;
 wire \channels.accum[2][13] ;
 wire \channels.accum[2][14] ;
 wire \channels.accum[2][15] ;
 wire \channels.accum[2][16] ;
 wire \channels.accum[2][17] ;
 wire \channels.accum[2][18] ;
 wire \channels.accum[2][19] ;
 wire \channels.accum[2][1] ;
 wire \channels.accum[2][20] ;
 wire \channels.accum[2][21] ;
 wire \channels.accum[2][22] ;
 wire \channels.accum[2][23] ;
 wire \channels.accum[2][2] ;
 wire \channels.accum[2][3] ;
 wire \channels.accum[2][4] ;
 wire \channels.accum[2][5] ;
 wire \channels.accum[2][6] ;
 wire \channels.accum[2][7] ;
 wire \channels.accum[2][8] ;
 wire \channels.accum[2][9] ;
 wire \channels.accum[3][0] ;
 wire \channels.accum[3][10] ;
 wire \channels.accum[3][11] ;
 wire \channels.accum[3][12] ;
 wire \channels.accum[3][13] ;
 wire \channels.accum[3][14] ;
 wire \channels.accum[3][15] ;
 wire \channels.accum[3][16] ;
 wire \channels.accum[3][17] ;
 wire \channels.accum[3][18] ;
 wire \channels.accum[3][19] ;
 wire \channels.accum[3][1] ;
 wire \channels.accum[3][20] ;
 wire \channels.accum[3][21] ;
 wire \channels.accum[3][22] ;
 wire \channels.accum[3][23] ;
 wire \channels.accum[3][2] ;
 wire \channels.accum[3][3] ;
 wire \channels.accum[3][4] ;
 wire \channels.accum[3][5] ;
 wire \channels.accum[3][6] ;
 wire \channels.accum[3][7] ;
 wire \channels.accum[3][8] ;
 wire \channels.accum[3][9] ;
 wire \channels.adsr_state[0][0] ;
 wire \channels.adsr_state[0][1] ;
 wire \channels.adsr_state[1][0] ;
 wire \channels.adsr_state[1][1] ;
 wire \channels.adsr_state[2][0] ;
 wire \channels.adsr_state[2][1] ;
 wire \channels.adsr_state[3][0] ;
 wire \channels.adsr_state[3][1] ;
 wire \channels.atk_dec1[0] ;
 wire \channels.atk_dec1[1] ;
 wire \channels.atk_dec1[2] ;
 wire \channels.atk_dec1[3] ;
 wire \channels.atk_dec1[4] ;
 wire \channels.atk_dec1[5] ;
 wire \channels.atk_dec1[6] ;
 wire \channels.atk_dec1[7] ;
 wire \channels.atk_dec2[0] ;
 wire \channels.atk_dec2[1] ;
 wire \channels.atk_dec2[2] ;
 wire \channels.atk_dec2[3] ;
 wire \channels.atk_dec2[4] ;
 wire \channels.atk_dec2[5] ;
 wire \channels.atk_dec2[6] ;
 wire \channels.atk_dec2[7] ;
 wire \channels.atk_dec3[0] ;
 wire \channels.atk_dec3[1] ;
 wire \channels.atk_dec3[2] ;
 wire \channels.atk_dec3[3] ;
 wire \channels.atk_dec3[4] ;
 wire \channels.atk_dec3[5] ;
 wire \channels.atk_dec3[6] ;
 wire \channels.atk_dec3[7] ;
 wire \channels.ch3_env[0] ;
 wire \channels.ch3_env[1] ;
 wire \channels.ch3_env[2] ;
 wire \channels.ch3_env[3] ;
 wire \channels.ch3_env[4] ;
 wire \channels.ch3_env[5] ;
 wire \channels.ch3_env[6] ;
 wire \channels.ch3_env[7] ;
 wire \channels.clk_div[0] ;
 wire \channels.clk_div[1] ;
 wire \channels.clk_div[2] ;
 wire \channels.ctrl_reg1[0] ;
 wire \channels.ctrl_reg1[1] ;
 wire \channels.ctrl_reg1[2] ;
 wire \channels.ctrl_reg1[3] ;
 wire \channels.ctrl_reg1[4] ;
 wire \channels.ctrl_reg1[5] ;
 wire \channels.ctrl_reg1[6] ;
 wire \channels.ctrl_reg1[7] ;
 wire \channels.ctrl_reg2[0] ;
 wire \channels.ctrl_reg2[1] ;
 wire \channels.ctrl_reg2[2] ;
 wire \channels.ctrl_reg2[3] ;
 wire \channels.ctrl_reg2[4] ;
 wire \channels.ctrl_reg2[5] ;
 wire \channels.ctrl_reg2[6] ;
 wire \channels.ctrl_reg2[7] ;
 wire \channels.ctrl_reg3[0] ;
 wire \channels.ctrl_reg3[1] ;
 wire \channels.ctrl_reg3[2] ;
 wire \channels.ctrl_reg3[3] ;
 wire \channels.ctrl_reg3[4] ;
 wire \channels.ctrl_reg3[5] ;
 wire \channels.ctrl_reg3[6] ;
 wire \channels.ctrl_reg3[7] ;
 wire \channels.env_counter[0][0] ;
 wire \channels.env_counter[0][10] ;
 wire \channels.env_counter[0][11] ;
 wire \channels.env_counter[0][12] ;
 wire \channels.env_counter[0][13] ;
 wire \channels.env_counter[0][14] ;
 wire \channels.env_counter[0][1] ;
 wire \channels.env_counter[0][2] ;
 wire \channels.env_counter[0][3] ;
 wire \channels.env_counter[0][4] ;
 wire \channels.env_counter[0][5] ;
 wire \channels.env_counter[0][6] ;
 wire \channels.env_counter[0][7] ;
 wire \channels.env_counter[0][8] ;
 wire \channels.env_counter[0][9] ;
 wire \channels.env_counter[1][0] ;
 wire \channels.env_counter[1][10] ;
 wire \channels.env_counter[1][11] ;
 wire \channels.env_counter[1][12] ;
 wire \channels.env_counter[1][13] ;
 wire \channels.env_counter[1][14] ;
 wire \channels.env_counter[1][1] ;
 wire \channels.env_counter[1][2] ;
 wire \channels.env_counter[1][3] ;
 wire \channels.env_counter[1][4] ;
 wire \channels.env_counter[1][5] ;
 wire \channels.env_counter[1][6] ;
 wire \channels.env_counter[1][7] ;
 wire \channels.env_counter[1][8] ;
 wire \channels.env_counter[1][9] ;
 wire \channels.env_counter[2][0] ;
 wire \channels.env_counter[2][10] ;
 wire \channels.env_counter[2][11] ;
 wire \channels.env_counter[2][12] ;
 wire \channels.env_counter[2][13] ;
 wire \channels.env_counter[2][14] ;
 wire \channels.env_counter[2][1] ;
 wire \channels.env_counter[2][2] ;
 wire \channels.env_counter[2][3] ;
 wire \channels.env_counter[2][4] ;
 wire \channels.env_counter[2][5] ;
 wire \channels.env_counter[2][6] ;
 wire \channels.env_counter[2][7] ;
 wire \channels.env_counter[2][8] ;
 wire \channels.env_counter[2][9] ;
 wire \channels.env_counter[3][0] ;
 wire \channels.env_counter[3][10] ;
 wire \channels.env_counter[3][11] ;
 wire \channels.env_counter[3][12] ;
 wire \channels.env_counter[3][13] ;
 wire \channels.env_counter[3][14] ;
 wire \channels.env_counter[3][1] ;
 wire \channels.env_counter[3][2] ;
 wire \channels.env_counter[3][3] ;
 wire \channels.env_counter[3][4] ;
 wire \channels.env_counter[3][5] ;
 wire \channels.env_counter[3][6] ;
 wire \channels.env_counter[3][7] ;
 wire \channels.env_counter[3][8] ;
 wire \channels.env_counter[3][9] ;
 wire \channels.env_vol[0][0] ;
 wire \channels.env_vol[0][1] ;
 wire \channels.env_vol[0][2] ;
 wire \channels.env_vol[0][3] ;
 wire \channels.env_vol[0][4] ;
 wire \channels.env_vol[0][5] ;
 wire \channels.env_vol[0][6] ;
 wire \channels.env_vol[0][7] ;
 wire \channels.env_vol[1][0] ;
 wire \channels.env_vol[1][1] ;
 wire \channels.env_vol[1][2] ;
 wire \channels.env_vol[1][3] ;
 wire \channels.env_vol[1][4] ;
 wire \channels.env_vol[1][5] ;
 wire \channels.env_vol[1][6] ;
 wire \channels.env_vol[1][7] ;
 wire \channels.env_vol[3][0] ;
 wire \channels.env_vol[3][1] ;
 wire \channels.env_vol[3][2] ;
 wire \channels.env_vol[3][3] ;
 wire \channels.env_vol[3][4] ;
 wire \channels.env_vol[3][5] ;
 wire \channels.env_vol[3][6] ;
 wire \channels.env_vol[3][7] ;
 wire \channels.exp_counter[0][0] ;
 wire \channels.exp_counter[0][1] ;
 wire \channels.exp_counter[0][2] ;
 wire \channels.exp_counter[0][3] ;
 wire \channels.exp_counter[0][4] ;
 wire \channels.exp_counter[1][0] ;
 wire \channels.exp_counter[1][1] ;
 wire \channels.exp_counter[1][2] ;
 wire \channels.exp_counter[1][3] ;
 wire \channels.exp_counter[1][4] ;
 wire \channels.exp_counter[2][0] ;
 wire \channels.exp_counter[2][1] ;
 wire \channels.exp_counter[2][2] ;
 wire \channels.exp_counter[2][3] ;
 wire \channels.exp_counter[2][4] ;
 wire \channels.exp_counter[3][0] ;
 wire \channels.exp_counter[3][1] ;
 wire \channels.exp_counter[3][2] ;
 wire \channels.exp_counter[3][3] ;
 wire \channels.exp_counter[3][4] ;
 wire \channels.exp_periods[0][0] ;
 wire \channels.exp_periods[0][1] ;
 wire \channels.exp_periods[0][2] ;
 wire \channels.exp_periods[0][3] ;
 wire \channels.exp_periods[0][4] ;
 wire \channels.exp_periods[1][0] ;
 wire \channels.exp_periods[1][1] ;
 wire \channels.exp_periods[1][2] ;
 wire \channels.exp_periods[1][3] ;
 wire \channels.exp_periods[1][4] ;
 wire \channels.exp_periods[2][0] ;
 wire \channels.exp_periods[2][1] ;
 wire \channels.exp_periods[2][2] ;
 wire \channels.exp_periods[2][3] ;
 wire \channels.exp_periods[2][4] ;
 wire \channels.exp_periods[3][0] ;
 wire \channels.exp_periods[3][1] ;
 wire \channels.exp_periods[3][2] ;
 wire \channels.exp_periods[3][3] ;
 wire \channels.exp_periods[3][4] ;
 wire \channels.freq1[0] ;
 wire \channels.freq1[10] ;
 wire \channels.freq1[11] ;
 wire \channels.freq1[12] ;
 wire \channels.freq1[13] ;
 wire \channels.freq1[14] ;
 wire \channels.freq1[15] ;
 wire \channels.freq1[1] ;
 wire \channels.freq1[2] ;
 wire \channels.freq1[3] ;
 wire \channels.freq1[4] ;
 wire \channels.freq1[5] ;
 wire \channels.freq1[6] ;
 wire \channels.freq1[7] ;
 wire \channels.freq1[8] ;
 wire \channels.freq1[9] ;
 wire \channels.freq2[0] ;
 wire \channels.freq2[10] ;
 wire \channels.freq2[11] ;
 wire \channels.freq2[12] ;
 wire \channels.freq2[13] ;
 wire \channels.freq2[14] ;
 wire \channels.freq2[15] ;
 wire \channels.freq2[1] ;
 wire \channels.freq2[2] ;
 wire \channels.freq2[3] ;
 wire \channels.freq2[4] ;
 wire \channels.freq2[5] ;
 wire \channels.freq2[6] ;
 wire \channels.freq2[7] ;
 wire \channels.freq2[8] ;
 wire \channels.freq2[9] ;
 wire \channels.freq3[0] ;
 wire \channels.freq3[10] ;
 wire \channels.freq3[11] ;
 wire \channels.freq3[12] ;
 wire \channels.freq3[13] ;
 wire \channels.freq3[14] ;
 wire \channels.freq3[15] ;
 wire \channels.freq3[1] ;
 wire \channels.freq3[2] ;
 wire \channels.freq3[3] ;
 wire \channels.freq3[4] ;
 wire \channels.freq3[5] ;
 wire \channels.freq3[6] ;
 wire \channels.freq3[7] ;
 wire \channels.freq3[8] ;
 wire \channels.freq3[9] ;
 wire \channels.lfsr[0][0] ;
 wire \channels.lfsr[0][10] ;
 wire \channels.lfsr[0][11] ;
 wire \channels.lfsr[0][12] ;
 wire \channels.lfsr[0][13] ;
 wire \channels.lfsr[0][14] ;
 wire \channels.lfsr[0][15] ;
 wire \channels.lfsr[0][16] ;
 wire \channels.lfsr[0][17] ;
 wire \channels.lfsr[0][18] ;
 wire \channels.lfsr[0][19] ;
 wire \channels.lfsr[0][1] ;
 wire \channels.lfsr[0][20] ;
 wire \channels.lfsr[0][21] ;
 wire \channels.lfsr[0][22] ;
 wire \channels.lfsr[0][2] ;
 wire \channels.lfsr[0][3] ;
 wire \channels.lfsr[0][4] ;
 wire \channels.lfsr[0][5] ;
 wire \channels.lfsr[0][6] ;
 wire \channels.lfsr[0][7] ;
 wire \channels.lfsr[0][8] ;
 wire \channels.lfsr[0][9] ;
 wire \channels.lfsr[1][0] ;
 wire \channels.lfsr[1][10] ;
 wire \channels.lfsr[1][11] ;
 wire \channels.lfsr[1][12] ;
 wire \channels.lfsr[1][13] ;
 wire \channels.lfsr[1][14] ;
 wire \channels.lfsr[1][15] ;
 wire \channels.lfsr[1][16] ;
 wire \channels.lfsr[1][17] ;
 wire \channels.lfsr[1][18] ;
 wire \channels.lfsr[1][19] ;
 wire \channels.lfsr[1][1] ;
 wire \channels.lfsr[1][20] ;
 wire \channels.lfsr[1][21] ;
 wire \channels.lfsr[1][22] ;
 wire \channels.lfsr[1][2] ;
 wire \channels.lfsr[1][3] ;
 wire \channels.lfsr[1][4] ;
 wire \channels.lfsr[1][5] ;
 wire \channels.lfsr[1][6] ;
 wire \channels.lfsr[1][7] ;
 wire \channels.lfsr[1][8] ;
 wire \channels.lfsr[1][9] ;
 wire \channels.lfsr[2][0] ;
 wire \channels.lfsr[2][10] ;
 wire \channels.lfsr[2][11] ;
 wire \channels.lfsr[2][12] ;
 wire \channels.lfsr[2][13] ;
 wire \channels.lfsr[2][14] ;
 wire \channels.lfsr[2][15] ;
 wire \channels.lfsr[2][16] ;
 wire \channels.lfsr[2][17] ;
 wire \channels.lfsr[2][18] ;
 wire \channels.lfsr[2][19] ;
 wire \channels.lfsr[2][1] ;
 wire \channels.lfsr[2][20] ;
 wire \channels.lfsr[2][21] ;
 wire \channels.lfsr[2][22] ;
 wire \channels.lfsr[2][2] ;
 wire \channels.lfsr[2][3] ;
 wire \channels.lfsr[2][4] ;
 wire \channels.lfsr[2][5] ;
 wire \channels.lfsr[2][6] ;
 wire \channels.lfsr[2][7] ;
 wire \channels.lfsr[2][8] ;
 wire \channels.lfsr[2][9] ;
 wire \channels.lfsr[3][0] ;
 wire \channels.lfsr[3][10] ;
 wire \channels.lfsr[3][11] ;
 wire \channels.lfsr[3][12] ;
 wire \channels.lfsr[3][13] ;
 wire \channels.lfsr[3][14] ;
 wire \channels.lfsr[3][15] ;
 wire \channels.lfsr[3][16] ;
 wire \channels.lfsr[3][17] ;
 wire \channels.lfsr[3][18] ;
 wire \channels.lfsr[3][19] ;
 wire \channels.lfsr[3][1] ;
 wire \channels.lfsr[3][20] ;
 wire \channels.lfsr[3][21] ;
 wire \channels.lfsr[3][22] ;
 wire \channels.lfsr[3][2] ;
 wire \channels.lfsr[3][3] ;
 wire \channels.lfsr[3][4] ;
 wire \channels.lfsr[3][5] ;
 wire \channels.lfsr[3][6] ;
 wire \channels.lfsr[3][7] ;
 wire \channels.lfsr[3][8] ;
 wire \channels.lfsr[3][9] ;
 wire \channels.pw1[0] ;
 wire \channels.pw1[10] ;
 wire \channels.pw1[11] ;
 wire \channels.pw1[1] ;
 wire \channels.pw1[2] ;
 wire \channels.pw1[3] ;
 wire \channels.pw1[4] ;
 wire \channels.pw1[5] ;
 wire \channels.pw1[6] ;
 wire \channels.pw1[7] ;
 wire \channels.pw1[8] ;
 wire \channels.pw1[9] ;
 wire \channels.pw2[0] ;
 wire \channels.pw2[10] ;
 wire \channels.pw2[11] ;
 wire \channels.pw2[1] ;
 wire \channels.pw2[2] ;
 wire \channels.pw2[3] ;
 wire \channels.pw2[4] ;
 wire \channels.pw2[5] ;
 wire \channels.pw2[6] ;
 wire \channels.pw2[7] ;
 wire \channels.pw2[8] ;
 wire \channels.pw2[9] ;
 wire \channels.pw3[0] ;
 wire \channels.pw3[10] ;
 wire \channels.pw3[11] ;
 wire \channels.pw3[1] ;
 wire \channels.pw3[2] ;
 wire \channels.pw3[3] ;
 wire \channels.pw3[4] ;
 wire \channels.pw3[5] ;
 wire \channels.pw3[6] ;
 wire \channels.pw3[7] ;
 wire \channels.pw3[8] ;
 wire \channels.pw3[9] ;
 wire \channels.ring_outs[0] ;
 wire \channels.ring_outs[1] ;
 wire \channels.ring_outs[2] ;
 wire \channels.sample1[0] ;
 wire \channels.sample1[10] ;
 wire \channels.sample1[11] ;
 wire \channels.sample1[1] ;
 wire \channels.sample1[2] ;
 wire \channels.sample1[3] ;
 wire \channels.sample1[4] ;
 wire \channels.sample1[5] ;
 wire \channels.sample1[6] ;
 wire \channels.sample1[7] ;
 wire \channels.sample1[8] ;
 wire \channels.sample1[9] ;
 wire \channels.sample2[0] ;
 wire \channels.sample2[10] ;
 wire \channels.sample2[11] ;
 wire \channels.sample2[1] ;
 wire \channels.sample2[2] ;
 wire \channels.sample2[3] ;
 wire \channels.sample2[4] ;
 wire \channels.sample2[5] ;
 wire \channels.sample2[6] ;
 wire \channels.sample2[7] ;
 wire \channels.sample2[8] ;
 wire \channels.sample2[9] ;
 wire \channels.sample3[0] ;
 wire \channels.sample3[10] ;
 wire \channels.sample3[11] ;
 wire \channels.sample3[1] ;
 wire \channels.sample3[2] ;
 wire \channels.sample3[3] ;
 wire \channels.sample3[4] ;
 wire \channels.sample3[5] ;
 wire \channels.sample3[6] ;
 wire \channels.sample3[7] ;
 wire \channels.sample3[8] ;
 wire \channels.sample3[9] ;
 wire \channels.sus_rel1[0] ;
 wire \channels.sus_rel1[1] ;
 wire \channels.sus_rel1[2] ;
 wire \channels.sus_rel1[3] ;
 wire \channels.sus_rel1[4] ;
 wire \channels.sus_rel1[5] ;
 wire \channels.sus_rel1[6] ;
 wire \channels.sus_rel1[7] ;
 wire \channels.sus_rel2[0] ;
 wire \channels.sus_rel2[1] ;
 wire \channels.sus_rel2[2] ;
 wire \channels.sus_rel2[3] ;
 wire \channels.sus_rel2[4] ;
 wire \channels.sus_rel2[5] ;
 wire \channels.sus_rel2[6] ;
 wire \channels.sus_rel2[7] ;
 wire \channels.sus_rel3[0] ;
 wire \channels.sus_rel3[1] ;
 wire \channels.sus_rel3[2] ;
 wire \channels.sus_rel3[3] ;
 wire \channels.sus_rel3[4] ;
 wire \channels.sus_rel3[5] ;
 wire \channels.sus_rel3[6] ;
 wire \channels.sus_rel3[7] ;
 wire \channels.sync_outs[0] ;
 wire \channels.sync_outs[1] ;
 wire \channels.sync_outs[2] ;
 wire \clk_ctr[0] ;
 wire \clk_ctr[1] ;
 wire \clk_trg[0] ;
 wire \clk_trg[1] ;
 wire clknet_0_clk;
 wire clknet_3_0_0_clk;
 wire clknet_3_1_0_clk;
 wire clknet_3_2_0_clk;
 wire clknet_3_3_0_clk;
 wire clknet_3_4_0_clk;
 wire clknet_3_5_0_clk;
 wire clknet_3_6_0_clk;
 wire clknet_3_7_0_clk;
 wire clknet_5_0__leaf_clk;
 wire clknet_5_10__leaf_clk;
 wire clknet_5_11__leaf_clk;
 wire clknet_5_12__leaf_clk;
 wire clknet_5_13__leaf_clk;
 wire clknet_5_14__leaf_clk;
 wire clknet_5_15__leaf_clk;
 wire clknet_5_16__leaf_clk;
 wire clknet_5_17__leaf_clk;
 wire clknet_5_18__leaf_clk;
 wire clknet_5_19__leaf_clk;
 wire clknet_5_1__leaf_clk;
 wire clknet_5_20__leaf_clk;
 wire clknet_5_21__leaf_clk;
 wire clknet_5_22__leaf_clk;
 wire clknet_5_23__leaf_clk;
 wire clknet_5_24__leaf_clk;
 wire clknet_5_25__leaf_clk;
 wire clknet_5_26__leaf_clk;
 wire clknet_5_27__leaf_clk;
 wire clknet_5_28__leaf_clk;
 wire clknet_5_29__leaf_clk;
 wire clknet_5_2__leaf_clk;
 wire clknet_5_30__leaf_clk;
 wire clknet_5_31__leaf_clk;
 wire clknet_5_3__leaf_clk;
 wire clknet_5_4__leaf_clk;
 wire clknet_5_5__leaf_clk;
 wire clknet_5_6__leaf_clk;
 wire clknet_5_7__leaf_clk;
 wire clknet_5_8__leaf_clk;
 wire clknet_5_9__leaf_clk;
 wire clknet_leaf_0_clk;
 wire clknet_leaf_100_clk;
 wire clknet_leaf_101_clk;
 wire clknet_leaf_102_clk;
 wire clknet_leaf_103_clk;
 wire clknet_leaf_104_clk;
 wire clknet_leaf_105_clk;
 wire clknet_leaf_106_clk;
 wire clknet_leaf_107_clk;
 wire clknet_leaf_108_clk;
 wire clknet_leaf_109_clk;
 wire clknet_leaf_110_clk;
 wire clknet_leaf_111_clk;
 wire clknet_leaf_112_clk;
 wire clknet_leaf_113_clk;
 wire clknet_leaf_114_clk;
 wire clknet_leaf_115_clk;
 wire clknet_leaf_116_clk;
 wire clknet_leaf_117_clk;
 wire clknet_leaf_118_clk;
 wire clknet_leaf_119_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_121_clk;
 wire clknet_leaf_122_clk;
 wire clknet_leaf_123_clk;
 wire clknet_leaf_124_clk;
 wire clknet_leaf_125_clk;
 wire clknet_leaf_127_clk;
 wire clknet_leaf_128_clk;
 wire clknet_leaf_129_clk;
 wire clknet_leaf_130_clk;
 wire clknet_leaf_131_clk;
 wire clknet_leaf_132_clk;
 wire clknet_leaf_133_clk;
 wire clknet_leaf_134_clk;
 wire clknet_leaf_135_clk;
 wire clknet_leaf_136_clk;
 wire clknet_leaf_137_clk;
 wire clknet_leaf_138_clk;
 wire clknet_leaf_139_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_141_clk;
 wire clknet_leaf_142_clk;
 wire clknet_leaf_143_clk;
 wire clknet_leaf_144_clk;
 wire clknet_leaf_145_clk;
 wire clknet_leaf_146_clk;
 wire clknet_leaf_147_clk;
 wire clknet_leaf_148_clk;
 wire clknet_leaf_149_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_150_clk;
 wire clknet_leaf_151_clk;
 wire clknet_leaf_152_clk;
 wire clknet_leaf_153_clk;
 wire clknet_leaf_154_clk;
 wire clknet_leaf_155_clk;
 wire clknet_leaf_156_clk;
 wire clknet_leaf_157_clk;
 wire clknet_leaf_158_clk;
 wire clknet_leaf_159_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_161_clk;
 wire clknet_leaf_162_clk;
 wire clknet_leaf_163_clk;
 wire clknet_leaf_164_clk;
 wire clknet_leaf_165_clk;
 wire clknet_leaf_166_clk;
 wire clknet_leaf_168_clk;
 wire clknet_leaf_169_clk;
 wire clknet_leaf_170_clk;
 wire clknet_leaf_171_clk;
 wire clknet_leaf_172_clk;
 wire clknet_leaf_173_clk;
 wire clknet_leaf_174_clk;
 wire clknet_leaf_175_clk;
 wire clknet_leaf_176_clk;
 wire clknet_leaf_177_clk;
 wire clknet_leaf_178_clk;
 wire clknet_leaf_179_clk;
 wire clknet_leaf_180_clk;
 wire clknet_leaf_181_clk;
 wire clknet_leaf_182_clk;
 wire clknet_leaf_185_clk;
 wire clknet_leaf_186_clk;
 wire clknet_leaf_187_clk;
 wire clknet_leaf_188_clk;
 wire clknet_leaf_189_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_190_clk;
 wire clknet_leaf_191_clk;
 wire clknet_leaf_192_clk;
 wire clknet_leaf_193_clk;
 wire clknet_leaf_194_clk;
 wire clknet_leaf_195_clk;
 wire clknet_leaf_196_clk;
 wire clknet_leaf_197_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_200_clk;
 wire clknet_leaf_201_clk;
 wire clknet_leaf_202_clk;
 wire clknet_leaf_203_clk;
 wire clknet_leaf_204_clk;
 wire clknet_leaf_205_clk;
 wire clknet_leaf_206_clk;
 wire clknet_leaf_207_clk;
 wire clknet_leaf_208_clk;
 wire clknet_leaf_209_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_210_clk;
 wire clknet_leaf_211_clk;
 wire clknet_leaf_212_clk;
 wire clknet_leaf_213_clk;
 wire clknet_leaf_214_clk;
 wire clknet_leaf_215_clk;
 wire clknet_leaf_216_clk;
 wire clknet_leaf_217_clk;
 wire clknet_leaf_218_clk;
 wire clknet_leaf_219_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_220_clk;
 wire clknet_leaf_221_clk;
 wire clknet_leaf_222_clk;
 wire clknet_leaf_223_clk;
 wire clknet_leaf_224_clk;
 wire clknet_leaf_225_clk;
 wire clknet_leaf_226_clk;
 wire clknet_leaf_227_clk;
 wire clknet_leaf_228_clk;
 wire clknet_leaf_229_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_230_clk;
 wire clknet_leaf_231_clk;
 wire clknet_leaf_232_clk;
 wire clknet_leaf_233_clk;
 wire clknet_leaf_235_clk;
 wire clknet_leaf_236_clk;
 wire clknet_leaf_238_clk;
 wire clknet_leaf_239_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_240_clk;
 wire clknet_leaf_242_clk;
 wire clknet_leaf_243_clk;
 wire clknet_leaf_244_clk;
 wire clknet_leaf_245_clk;
 wire clknet_leaf_246_clk;
 wire clknet_leaf_247_clk;
 wire clknet_leaf_248_clk;
 wire clknet_leaf_249_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_52_clk;
 wire clknet_leaf_53_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_55_clk;
 wire clknet_leaf_56_clk;
 wire clknet_leaf_57_clk;
 wire clknet_leaf_58_clk;
 wire clknet_leaf_59_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_60_clk;
 wire clknet_leaf_61_clk;
 wire clknet_leaf_62_clk;
 wire clknet_leaf_63_clk;
 wire clknet_leaf_64_clk;
 wire clknet_leaf_66_clk;
 wire clknet_leaf_67_clk;
 wire clknet_leaf_68_clk;
 wire clknet_leaf_69_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_70_clk;
 wire clknet_leaf_71_clk;
 wire clknet_leaf_72_clk;
 wire clknet_leaf_73_clk;
 wire clknet_leaf_74_clk;
 wire clknet_leaf_75_clk;
 wire clknet_leaf_76_clk;
 wire clknet_leaf_77_clk;
 wire clknet_leaf_78_clk;
 wire clknet_leaf_79_clk;
 wire clknet_leaf_80_clk;
 wire clknet_leaf_81_clk;
 wire clknet_leaf_82_clk;
 wire clknet_leaf_85_clk;
 wire clknet_leaf_86_clk;
 wire clknet_leaf_87_clk;
 wire clknet_leaf_88_clk;
 wire clknet_leaf_89_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_90_clk;
 wire clknet_leaf_91_clk;
 wire clknet_leaf_93_clk;
 wire clknet_leaf_94_clk;
 wire clknet_leaf_95_clk;
 wire clknet_leaf_96_clk;
 wire clknet_leaf_97_clk;
 wire clknet_leaf_98_clk;
 wire clknet_leaf_99_clk;
 wire clknet_leaf_9_clk;
 wire \filters.band[0] ;
 wire \filters.band[10] ;
 wire \filters.band[11] ;
 wire \filters.band[12] ;
 wire \filters.band[13] ;
 wire \filters.band[14] ;
 wire \filters.band[15] ;
 wire \filters.band[16] ;
 wire \filters.band[17] ;
 wire \filters.band[18] ;
 wire \filters.band[19] ;
 wire \filters.band[1] ;
 wire \filters.band[20] ;
 wire \filters.band[21] ;
 wire \filters.band[22] ;
 wire \filters.band[23] ;
 wire \filters.band[24] ;
 wire \filters.band[25] ;
 wire \filters.band[26] ;
 wire \filters.band[27] ;
 wire \filters.band[28] ;
 wire \filters.band[29] ;
 wire \filters.band[2] ;
 wire \filters.band[30] ;
 wire \filters.band[31] ;
 wire \filters.band[3] ;
 wire \filters.band[4] ;
 wire \filters.band[5] ;
 wire \filters.band[6] ;
 wire \filters.band[7] ;
 wire \filters.band[8] ;
 wire \filters.band[9] ;
 wire \filters.bp ;
 wire \filters.cutoff_lut[10] ;
 wire \filters.cutoff_lut[11] ;
 wire \filters.cutoff_lut[12] ;
 wire \filters.cutoff_lut[13] ;
 wire \filters.cutoff_lut[14] ;
 wire \filters.cutoff_lut[15] ;
 wire \filters.cutoff_lut[16] ;
 wire \filters.cutoff_lut[6] ;
 wire \filters.cutoff_lut[7] ;
 wire \filters.cutoff_lut[8] ;
 wire \filters.cutoff_lut[9] ;
 wire \filters.filt_1 ;
 wire \filters.filt_2 ;
 wire \filters.filt_3 ;
 wire \filters.filter_step[0] ;
 wire \filters.filter_step[1] ;
 wire \filters.filter_step[2] ;
 wire \filters.high[0] ;
 wire \filters.high[10] ;
 wire \filters.high[11] ;
 wire \filters.high[12] ;
 wire \filters.high[13] ;
 wire \filters.high[14] ;
 wire \filters.high[15] ;
 wire \filters.high[16] ;
 wire \filters.high[17] ;
 wire \filters.high[18] ;
 wire \filters.high[19] ;
 wire \filters.high[1] ;
 wire \filters.high[20] ;
 wire \filters.high[21] ;
 wire \filters.high[22] ;
 wire \filters.high[23] ;
 wire \filters.high[24] ;
 wire \filters.high[25] ;
 wire \filters.high[26] ;
 wire \filters.high[27] ;
 wire \filters.high[28] ;
 wire \filters.high[29] ;
 wire \filters.high[2] ;
 wire \filters.high[30] ;
 wire \filters.high[31] ;
 wire \filters.high[3] ;
 wire \filters.high[4] ;
 wire \filters.high[5] ;
 wire \filters.high[6] ;
 wire \filters.high[7] ;
 wire \filters.high[8] ;
 wire \filters.high[9] ;
 wire \filters.hp ;
 wire \filters.low[0] ;
 wire \filters.low[10] ;
 wire \filters.low[11] ;
 wire \filters.low[12] ;
 wire \filters.low[13] ;
 wire \filters.low[14] ;
 wire \filters.low[15] ;
 wire \filters.low[16] ;
 wire \filters.low[17] ;
 wire \filters.low[18] ;
 wire \filters.low[19] ;
 wire \filters.low[1] ;
 wire \filters.low[20] ;
 wire \filters.low[21] ;
 wire \filters.low[22] ;
 wire \filters.low[23] ;
 wire \filters.low[24] ;
 wire \filters.low[25] ;
 wire \filters.low[26] ;
 wire \filters.low[27] ;
 wire \filters.low[28] ;
 wire \filters.low[29] ;
 wire \filters.low[2] ;
 wire \filters.low[30] ;
 wire \filters.low[31] ;
 wire \filters.low[3] ;
 wire \filters.low[4] ;
 wire \filters.low[5] ;
 wire \filters.low[6] ;
 wire \filters.low[7] ;
 wire \filters.low[8] ;
 wire \filters.low[9] ;
 wire \filters.lp ;
 wire \filters.mode_vol[0] ;
 wire \filters.mode_vol[1] ;
 wire \filters.mode_vol[2] ;
 wire \filters.mode_vol[3] ;
 wire \filters.mode_vol[7] ;
 wire \filters.res_filt[3] ;
 wire \filters.res_filt[4] ;
 wire \filters.res_filt[5] ;
 wire \filters.res_filt[6] ;
 wire \filters.res_filt[7] ;
 wire \filters.res_lut[0] ;
 wire \filters.res_lut[10] ;
 wire \filters.res_lut[1] ;
 wire \filters.res_lut[2] ;
 wire \filters.res_lut[3] ;
 wire \filters.res_lut[4] ;
 wire \filters.res_lut[5] ;
 wire \filters.res_lut[6] ;
 wire \filters.res_lut[7] ;
 wire \filters.res_lut[8] ;
 wire \filters.res_lut[9] ;
 wire \filters.sample_buff[0] ;
 wire \filters.sample_buff[10] ;
 wire \filters.sample_buff[11] ;
 wire \filters.sample_buff[12] ;
 wire \filters.sample_buff[13] ;
 wire \filters.sample_buff[14] ;
 wire \filters.sample_buff[1] ;
 wire \filters.sample_buff[2] ;
 wire \filters.sample_buff[3] ;
 wire \filters.sample_buff[4] ;
 wire \filters.sample_buff[5] ;
 wire \filters.sample_buff[6] ;
 wire \filters.sample_buff[7] ;
 wire \filters.sample_buff[8] ;
 wire \filters.sample_buff[9] ;
 wire \filters.sample_filtered[0] ;
 wire \filters.sample_filtered[10] ;
 wire \filters.sample_filtered[11] ;
 wire \filters.sample_filtered[12] ;
 wire \filters.sample_filtered[13] ;
 wire \filters.sample_filtered[14] ;
 wire \filters.sample_filtered[15] ;
 wire \filters.sample_filtered[1] ;
 wire \filters.sample_filtered[2] ;
 wire \filters.sample_filtered[3] ;
 wire \filters.sample_filtered[4] ;
 wire \filters.sample_filtered[5] ;
 wire \filters.sample_filtered[6] ;
 wire \filters.sample_filtered[7] ;
 wire \filters.sample_filtered[8] ;
 wire \filters.sample_filtered[9] ;
 wire net1;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net2;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net3;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net4;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net5;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net6;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net8;
 wire net9;
 wire \spi_dac_i.counter[0] ;
 wire \spi_dac_i.counter[1] ;
 wire \spi_dac_i.counter[2] ;
 wire \spi_dac_i.counter[3] ;
 wire \spi_dac_i.counter[4] ;
 wire \spi_dac_i.spi_dat_buff_0[0] ;
 wire \spi_dac_i.spi_dat_buff_0[10] ;
 wire \spi_dac_i.spi_dat_buff_0[11] ;
 wire \spi_dac_i.spi_dat_buff_0[1] ;
 wire \spi_dac_i.spi_dat_buff_0[2] ;
 wire \spi_dac_i.spi_dat_buff_0[3] ;
 wire \spi_dac_i.spi_dat_buff_0[4] ;
 wire \spi_dac_i.spi_dat_buff_0[5] ;
 wire \spi_dac_i.spi_dat_buff_0[6] ;
 wire \spi_dac_i.spi_dat_buff_0[7] ;
 wire \spi_dac_i.spi_dat_buff_0[8] ;
 wire \spi_dac_i.spi_dat_buff_0[9] ;
 wire \spi_dac_i.spi_dat_buff_1[0] ;
 wire \spi_dac_i.spi_dat_buff_1[10] ;
 wire \spi_dac_i.spi_dat_buff_1[11] ;
 wire \spi_dac_i.spi_dat_buff_1[1] ;
 wire \spi_dac_i.spi_dat_buff_1[2] ;
 wire \spi_dac_i.spi_dat_buff_1[3] ;
 wire \spi_dac_i.spi_dat_buff_1[4] ;
 wire \spi_dac_i.spi_dat_buff_1[5] ;
 wire \spi_dac_i.spi_dat_buff_1[6] ;
 wire \spi_dac_i.spi_dat_buff_1[7] ;
 wire \spi_dac_i.spi_dat_buff_1[8] ;
 wire \spi_dac_i.spi_dat_buff_1[9] ;
 wire \tt_um_rejunity_sn76489.chan[0].attenuation.control[0] ;
 wire \tt_um_rejunity_sn76489.chan[0].attenuation.control[1] ;
 wire \tt_um_rejunity_sn76489.chan[0].attenuation.control[2] ;
 wire \tt_um_rejunity_sn76489.chan[0].attenuation.control[3] ;
 wire \tt_um_rejunity_sn76489.chan[0].attenuation.in ;
 wire \tt_um_rejunity_sn76489.chan[1].attenuation.control[0] ;
 wire \tt_um_rejunity_sn76489.chan[1].attenuation.control[1] ;
 wire \tt_um_rejunity_sn76489.chan[1].attenuation.control[2] ;
 wire \tt_um_rejunity_sn76489.chan[1].attenuation.control[3] ;
 wire \tt_um_rejunity_sn76489.chan[1].attenuation.in ;
 wire \tt_um_rejunity_sn76489.chan[2].attenuation.control[0] ;
 wire \tt_um_rejunity_sn76489.chan[2].attenuation.control[1] ;
 wire \tt_um_rejunity_sn76489.chan[2].attenuation.control[2] ;
 wire \tt_um_rejunity_sn76489.chan[2].attenuation.control[3] ;
 wire \tt_um_rejunity_sn76489.chan[2].attenuation.in ;
 wire \tt_um_rejunity_sn76489.chan[3].attenuation.control[0] ;
 wire \tt_um_rejunity_sn76489.chan[3].attenuation.control[1] ;
 wire \tt_um_rejunity_sn76489.chan[3].attenuation.control[2] ;
 wire \tt_um_rejunity_sn76489.chan[3].attenuation.control[3] ;
 wire \tt_um_rejunity_sn76489.chan[3].attenuation.in ;
 wire \tt_um_rejunity_sn76489.clk_counter[0] ;
 wire \tt_um_rejunity_sn76489.clk_counter[1] ;
 wire \tt_um_rejunity_sn76489.clk_counter[2] ;
 wire \tt_um_rejunity_sn76489.clk_counter[3] ;
 wire \tt_um_rejunity_sn76489.clk_counter[4] ;
 wire \tt_um_rejunity_sn76489.control_noise[0][0] ;
 wire \tt_um_rejunity_sn76489.control_noise[0][1] ;
 wire \tt_um_rejunity_sn76489.control_noise[0][2] ;
 wire \tt_um_rejunity_sn76489.control_tone_freq[0][0] ;
 wire \tt_um_rejunity_sn76489.control_tone_freq[0][1] ;
 wire \tt_um_rejunity_sn76489.control_tone_freq[0][2] ;
 wire \tt_um_rejunity_sn76489.control_tone_freq[0][3] ;
 wire \tt_um_rejunity_sn76489.control_tone_freq[0][4] ;
 wire \tt_um_rejunity_sn76489.control_tone_freq[0][5] ;
 wire \tt_um_rejunity_sn76489.control_tone_freq[0][6] ;
 wire \tt_um_rejunity_sn76489.control_tone_freq[0][7] ;
 wire \tt_um_rejunity_sn76489.control_tone_freq[0][8] ;
 wire \tt_um_rejunity_sn76489.control_tone_freq[0][9] ;
 wire \tt_um_rejunity_sn76489.control_tone_freq[1][0] ;
 wire \tt_um_rejunity_sn76489.control_tone_freq[1][1] ;
 wire \tt_um_rejunity_sn76489.control_tone_freq[1][2] ;
 wire \tt_um_rejunity_sn76489.control_tone_freq[1][3] ;
 wire \tt_um_rejunity_sn76489.control_tone_freq[1][4] ;
 wire \tt_um_rejunity_sn76489.control_tone_freq[1][5] ;
 wire \tt_um_rejunity_sn76489.control_tone_freq[1][6] ;
 wire \tt_um_rejunity_sn76489.control_tone_freq[1][7] ;
 wire \tt_um_rejunity_sn76489.control_tone_freq[1][8] ;
 wire \tt_um_rejunity_sn76489.control_tone_freq[1][9] ;
 wire \tt_um_rejunity_sn76489.control_tone_freq[2][0] ;
 wire \tt_um_rejunity_sn76489.control_tone_freq[2][1] ;
 wire \tt_um_rejunity_sn76489.control_tone_freq[2][2] ;
 wire \tt_um_rejunity_sn76489.control_tone_freq[2][3] ;
 wire \tt_um_rejunity_sn76489.control_tone_freq[2][4] ;
 wire \tt_um_rejunity_sn76489.control_tone_freq[2][5] ;
 wire \tt_um_rejunity_sn76489.control_tone_freq[2][6] ;
 wire \tt_um_rejunity_sn76489.control_tone_freq[2][7] ;
 wire \tt_um_rejunity_sn76489.control_tone_freq[2][8] ;
 wire \tt_um_rejunity_sn76489.control_tone_freq[2][9] ;
 wire \tt_um_rejunity_sn76489.latch_control_reg[0] ;
 wire \tt_um_rejunity_sn76489.latch_control_reg[1] ;
 wire \tt_um_rejunity_sn76489.latch_control_reg[2] ;
 wire \tt_um_rejunity_sn76489.noise[0].gen.counter[0] ;
 wire \tt_um_rejunity_sn76489.noise[0].gen.counter[1] ;
 wire \tt_um_rejunity_sn76489.noise[0].gen.counter[2] ;
 wire \tt_um_rejunity_sn76489.noise[0].gen.counter[3] ;
 wire \tt_um_rejunity_sn76489.noise[0].gen.counter[4] ;
 wire \tt_um_rejunity_sn76489.noise[0].gen.counter[5] ;
 wire \tt_um_rejunity_sn76489.noise[0].gen.counter[6] ;
 wire \tt_um_rejunity_sn76489.noise[0].gen.lfsr[10] ;
 wire \tt_um_rejunity_sn76489.noise[0].gen.lfsr[11] ;
 wire \tt_um_rejunity_sn76489.noise[0].gen.lfsr[12] ;
 wire \tt_um_rejunity_sn76489.noise[0].gen.lfsr[13] ;
 wire \tt_um_rejunity_sn76489.noise[0].gen.lfsr[14] ;
 wire \tt_um_rejunity_sn76489.noise[0].gen.lfsr[1] ;
 wire \tt_um_rejunity_sn76489.noise[0].gen.lfsr[2] ;
 wire \tt_um_rejunity_sn76489.noise[0].gen.lfsr[3] ;
 wire \tt_um_rejunity_sn76489.noise[0].gen.lfsr[4] ;
 wire \tt_um_rejunity_sn76489.noise[0].gen.lfsr[5] ;
 wire \tt_um_rejunity_sn76489.noise[0].gen.lfsr[6] ;
 wire \tt_um_rejunity_sn76489.noise[0].gen.lfsr[7] ;
 wire \tt_um_rejunity_sn76489.noise[0].gen.lfsr[8] ;
 wire \tt_um_rejunity_sn76489.noise[0].gen.lfsr[9] ;
 wire \tt_um_rejunity_sn76489.noise[0].gen.restart_noise ;
 wire \tt_um_rejunity_sn76489.noise[0].gen.signal_edge.previous_signal_state_0 ;
 wire \tt_um_rejunity_sn76489.tone[0].gen.counter[0] ;
 wire \tt_um_rejunity_sn76489.tone[0].gen.counter[1] ;
 wire \tt_um_rejunity_sn76489.tone[0].gen.counter[2] ;
 wire \tt_um_rejunity_sn76489.tone[0].gen.counter[3] ;
 wire \tt_um_rejunity_sn76489.tone[0].gen.counter[4] ;
 wire \tt_um_rejunity_sn76489.tone[0].gen.counter[5] ;
 wire \tt_um_rejunity_sn76489.tone[0].gen.counter[6] ;
 wire \tt_um_rejunity_sn76489.tone[0].gen.counter[7] ;
 wire \tt_um_rejunity_sn76489.tone[0].gen.counter[8] ;
 wire \tt_um_rejunity_sn76489.tone[0].gen.counter[9] ;
 wire \tt_um_rejunity_sn76489.tone[1].gen.counter[0] ;
 wire \tt_um_rejunity_sn76489.tone[1].gen.counter[1] ;
 wire \tt_um_rejunity_sn76489.tone[1].gen.counter[2] ;
 wire \tt_um_rejunity_sn76489.tone[1].gen.counter[3] ;
 wire \tt_um_rejunity_sn76489.tone[1].gen.counter[4] ;
 wire \tt_um_rejunity_sn76489.tone[1].gen.counter[5] ;
 wire \tt_um_rejunity_sn76489.tone[1].gen.counter[6] ;
 wire \tt_um_rejunity_sn76489.tone[1].gen.counter[7] ;
 wire \tt_um_rejunity_sn76489.tone[1].gen.counter[8] ;
 wire \tt_um_rejunity_sn76489.tone[1].gen.counter[9] ;
 wire \tt_um_rejunity_sn76489.tone[2].gen.counter[0] ;
 wire \tt_um_rejunity_sn76489.tone[2].gen.counter[1] ;
 wire \tt_um_rejunity_sn76489.tone[2].gen.counter[2] ;
 wire \tt_um_rejunity_sn76489.tone[2].gen.counter[3] ;
 wire \tt_um_rejunity_sn76489.tone[2].gen.counter[4] ;
 wire \tt_um_rejunity_sn76489.tone[2].gen.counter[5] ;
 wire \tt_um_rejunity_sn76489.tone[2].gen.counter[6] ;
 wire \tt_um_rejunity_sn76489.tone[2].gen.counter[7] ;
 wire \tt_um_rejunity_sn76489.tone[2].gen.counter[8] ;
 wire \tt_um_rejunity_sn76489.tone[2].gen.counter[9] ;

 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_1 (.I(_01588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_10 (.I(_01590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_2 (.I(_01588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_3 (.I(_01590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_4 (.I(_01588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_5 (.I(_01590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_6 (.I(_01590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_7 (.I(_01590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_8 (.I(_01590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_9 (.I(_01590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08467__I (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08468__I (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08469__A1 (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08470__A2 (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08471__A1 (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08471__A2 (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08474__A2 (.I(_01003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08475__I (.I(_01004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08477__A1 (.I(_01006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08478__A1 (.I(\filters.res_filt[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08479__I (.I(_01008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08480__I (.I(net17));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08481__A2 (.I(_01003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08482__A1 (.I(net14));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08483__I (.I(_01004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08484__A1 (.I(\filters.res_filt[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08484__A2 (.I(_01013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08485__A2 (.I(_01012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08486__I (.I(_01015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08488__A1 (.I(_01017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08490__A2 (.I(_01019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08492__A2 (.I(_00129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08493__A1 (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08494__A1 (.I(\filters.res_filt[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08494__A2 (.I(_01013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08495__A2 (.I(_01022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08496__I (.I(_01024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08497__I (.I(_01015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08498__A2 (.I(_01019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08500__I (.I(_01024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08503__A2 (.I(_00129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08505__A1 (.I(_01008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08505__A2 (.I(_01019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08505__B (.I(_01032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08513__I (.I(_01008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08514__B (.I(_00129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08515__I (.I(net17));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08516__I (.I(_01042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08517__A1 (.I(_01043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08517__A2 (.I(_01008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08518__A1 (.I(_01024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08526__A1 (.I(_01043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08539__I0 (.I(_01019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08545__I (.I(net17));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08547__A1 (.I(\clk_trg[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08548__I (.I(\clk_trg[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08551__A1 (.I(\clk_trg[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08551__B2 (.I(\clk_trg[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08552__A1 (.I(_01062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08553__A1 (.I(\channels.clk_div[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08553__A2 (.I(_01069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08566__A1 (.I(_01070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08566__A2 (.I(_01082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08567__I (.I(_01083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08568__S0 (.I(_00009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08568__S1 (.I(_00010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08569__I (.I(_01085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08570__I (.I(_01042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08571__A2 (.I(_01083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08573__I (.I(_01089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08574__A2 (.I(_01086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08574__B1 (.I(_01090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08574__B2 (.I(\channels.ring_outs[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08576__I (.I(\channels.clk_div[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08578__A1 (.I(net17));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08578__A2 (.I(_01093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08584__A2 (.I(_01099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08585__I (.I(_01100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08586__I (.I(_01042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08587__A1 (.I(_01102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08587__A2 (.I(_01100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08589__I (.I(_01104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08590__A1 (.I(_01086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08590__B1 (.I(_01105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08590__B2 (.I(\channels.ring_outs[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08654__I (.I(_00009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08655__I (.I(_01138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08656__I (.I(_01139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08657__I (.I(_01140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08658__I (.I(_01141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08659__I (.I(_01142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08661__I (.I(_01144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08662__I (.I(_01145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08663__I (.I(_01146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08664__I (.I(_01147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08665__I (.I(_01148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08666__I (.I(_01149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08667__I (.I(_01150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08668__I (.I(_01151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08669__I (.I(_00010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08671__I (.I(_01154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08672__I (.I(_01155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08676__I (.I(_01159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08677__I (.I(_01160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08678__I (.I(_01161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08679__I (.I(_01162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08680__I (.I(_01163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08681__I (.I(_01164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08682__I (.I(_01165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08683__I (.I(_01166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08684__I (.I(_01167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08685__S0 (.I(_01152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08685__S1 (.I(_01168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08686__I (.I(_01165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08687__I (.I(_01170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08688__I (.I(_01171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08689__I (.I(_01172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08691__I (.I(_01152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08700__A1 (.I(_01169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08701__S1 (.I(_01172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08707__S1 (.I(_01172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08714__S1 (.I(_01172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08720__A1 (.I(_01201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08722__S0 (.I(_01152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08722__S1 (.I(_01168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08734__A1 (.I(_01169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08735__I (.I(_01100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08736__I (.I(_01219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08737__A2 (.I(_01105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08739__A1 (.I(_01169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08740__A1 (.I(_01169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08743__A2 (.I(_01105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08747__A2 (.I(_01105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08755__A2 (.I(_01230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08759__A2 (.I(_01230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08761__I (.I(_01083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08762__I (.I(_01240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08763__A2 (.I(_01090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08765__A2 (.I(_01090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08767__A2 (.I(_01090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08770__A2 (.I(_01245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08772__A2 (.I(_01245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08780__I (.I(_01253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08781__I (.I(_01254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08782__A1 (.I(_01102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08782__A2 (.I(_01253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08784__I (.I(_01257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08785__A1 (.I(_01086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08785__B1 (.I(_01258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08785__B2 (.I(\channels.ring_outs[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08789__I (.I(_01261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08795__A2 (.I(\channels.ctrl_reg2[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08796__A2 (.I(\channels.ctrl_reg3[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08796__B1 (.I(\channels.ctrl_reg1[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08798__A1 (.I(\channels.ctrl_reg3[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08798__A3 (.I(_01082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08810__A1 (.I(\channels.ctrl_reg2[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08810__A3 (.I(_01282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08814__I (.I(_01286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08823__A1 (.I(\channels.ctrl_reg1[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08823__A3 (.I(_01295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08825__A1 (.I(_01270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08828__A1 (.I(\channels.freq3[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08829__B2 (.I(\channels.freq1[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08832__I (.I(_01142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08833__I (.I(_01305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08835__I (.I(_01307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08836__A1 (.I(_01308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08837__A1 (.I(_01146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08839__A1 (.I(_01308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08840__A1 (.I(_01308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08840__C (.I(_01159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08841__A1 (.I(_01304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08842__A1 (.I(_01303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08843__A1 (.I(_01300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08844__I (.I(_01253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08845__I (.I(_01317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08847__I (.I(_01295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08848__A1 (.I(_01070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08848__A2 (.I(_01319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08849__I (.I(_01320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08850__I (.I(_01321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08852__A1 (.I(_01160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08852__C (.I(_01303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08853__A1 (.I(\channels.freq3[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08854__B2 (.I(\channels.freq1[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08857__S0 (.I(_01307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08857__S1 (.I(_01328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08858__A1 (.I(_01327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08861__A1 (.I(_01323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08863__A2 (.I(_01334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08867__A1 (.I(_01327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08868__A1 (.I(\channels.freq3[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08869__A1 (.I(\channels.freq2[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08869__B2 (.I(\channels.freq1[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08871__S0 (.I(_01145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08871__S1 (.I(_01159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08872__A1 (.I(_01341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08872__A2 (.I(_01342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08877__A1 (.I(_01337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08880__A1 (.I(_01341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08880__A2 (.I(_01342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08882__A1 (.I(\channels.freq3[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08883__B2 (.I(\channels.freq1[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08885__S0 (.I(_01308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08885__S1 (.I(_01160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08886__A1 (.I(_01354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08889__A1 (.I(_01349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08890__I (.I(_01257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08891__A2 (.I(_01360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08895__A1 (.I(_01354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08896__A1 (.I(\channels.freq3[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08897__B2 (.I(\channels.freq1[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08899__S0 (.I(_01146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08899__S1 (.I(_01161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08900__A1 (.I(_01367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08900__A2 (.I(_01368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08903__A1 (.I(_01337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08904__B1 (.I(_01372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08905__A1 (.I(_01367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08905__A2 (.I(_01368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08908__B2 (.I(\channels.freq1[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08910__S0 (.I(_01147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08910__S1 (.I(_01161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08911__A1 (.I(_01377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08913__A1 (.I(_01349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08914__A2 (.I(_01360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08917__A1 (.I(_01377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08921__B2 (.I(\channels.freq1[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08923__S0 (.I(_01147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08923__S1 (.I(_01162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08924__A1 (.I(_01389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08928__A1 (.I(_01337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08930__A1 (.I(_01389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08932__A1 (.I(\channels.freq3[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08933__B2 (.I(\channels.freq1[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08935__S0 (.I(_01148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08935__S1 (.I(_01163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08936__A1 (.I(_01400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08940__A1 (.I(_01349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08941__A2 (.I(_01360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08944__I (.I(_01257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08945__A1 (.I(_01400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08948__A1 (.I(\channels.freq2[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08948__B2 (.I(\channels.freq1[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08950__S0 (.I(_01148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08950__S1 (.I(_01163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08951__A1 (.I(_01414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08951__A2 (.I(_01415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08955__A1 (.I(_01337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08956__I (.I(_01254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08957__B1 (.I(_01420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08958__I (.I(_01321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08959__A1 (.I(_01414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08959__A2 (.I(_01415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08962__A1 (.I(\channels.freq2[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08962__B2 (.I(\channels.freq1[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08964__S0 (.I(_01148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08964__S1 (.I(_01163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08965__A1 (.I(_01427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08969__A1 (.I(_01349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08970__A2 (.I(_01360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08971__A1 (.I(_01422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08974__A1 (.I(_01427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08977__A1 (.I(\channels.freq3[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08978__A1 (.I(\channels.freq2[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08978__B2 (.I(\channels.freq1[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08980__S0 (.I(_01149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08980__S1 (.I(_01164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08981__A1 (.I(_01442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08981__A2 (.I(_01443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08985__A1 (.I(_01436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08986__B1 (.I(_01448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08988__A1 (.I(_01442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08988__A2 (.I(_01443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08990__A1 (.I(\channels.freq2[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08990__B2 (.I(\channels.freq1[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08992__S0 (.I(_01149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08992__S1 (.I(_01165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08993__A1 (.I(_01453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08997__A1 (.I(_01449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08999__I (.I(_01460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09000__A2 (.I(_01461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09001__A1 (.I(_01422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09003__A1 (.I(_01453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09006__A1 (.I(\channels.freq2[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09006__B2 (.I(\channels.freq1[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09008__S0 (.I(_01140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09008__S1 (.I(_01154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09009__I (.I(_01469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09010__A1 (.I(_01468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09010__A2 (.I(_01470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09014__A1 (.I(_01436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09015__B1 (.I(_01475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09016__A1 (.I(_01468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09016__A2 (.I(_01470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09018__A1 (.I(\channels.freq2[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09018__B2 (.I(\channels.freq1[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09020__I (.I(_00010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09021__S0 (.I(_01138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09021__S1 (.I(_01480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09022__I (.I(_01481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09023__A1 (.I(_01479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09023__A2 (.I(_01482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09027__A1 (.I(_01449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09028__A2 (.I(_01461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09029__A1 (.I(_01422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09031__A1 (.I(_01479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09031__A2 (.I(_01482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09034__A1 (.I(\channels.freq2[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09034__B2 (.I(\channels.freq1[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09036__I (.I(_01138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09038__S0 (.I(_01495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09038__S1 (.I(_01496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09039__I (.I(_01497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09040__A1 (.I(_01494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09044__A1 (.I(_01436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09045__B1 (.I(_01503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09046__A1 (.I(_01494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09046__A2 (.I(_01497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09048__A1 (.I(\channels.freq2[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09048__B2 (.I(\channels.freq1[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09049__A1 (.I(_01505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09049__A2 (.I(_01506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09050__S0 (.I(_00009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09051__I (.I(_01508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09053__A2 (.I(_01510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09057__A1 (.I(_01449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09058__A2 (.I(_01461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09059__A1 (.I(_01422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09061__I (.I(_01257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09062__A1 (.I(_01505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09062__A2 (.I(_01506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09062__B (.I(_01510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09063__S0 (.I(_01139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09063__S1 (.I(_01480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09064__I (.I(_01520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09065__A3 (.I(_01521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09066__B (.I(_01521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09067__A1 (.I(_01436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09068__I (.I(_01254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09069__B1 (.I(_01524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09071__S0 (.I(_01139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09071__S1 (.I(_01480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09072__I (.I(_01527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09073__A2 (.I(_01528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09074__A1 (.I(_01323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09075__A2 (.I(_01334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09075__B1 (.I(_01530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09078__S0 (.I(_01495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09078__S1 (.I(_01496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09079__I (.I(_01533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09080__A2 (.I(_01528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09080__B (.I(_01534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09081__A2 (.I(_01528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09081__A3 (.I(_01534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09083__A1 (.I(_01323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09085__B1 (.I(_01539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09086__I (.I(_01321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09087__S0 (.I(_01495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09087__S1 (.I(_01496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09088__I (.I(_01541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09089__I (.I(_01542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09091__A1 (.I(_01449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09092__A2 (.I(_01461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09093__A1 (.I(_01540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09096__S0 (.I(_01138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09097__I (.I(_01549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09098__A2 (.I(_01550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09099__A1 (.I(_01300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09100__B1 (.I(_01552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09101__I (.I(_01549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09103__S0 (.I(_01139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09103__S1 (.I(_01480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09104__I (.I(_01555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09105__A2 (.I(_01556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09106__A2 (.I(_01556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09107__A1 (.I(_01323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09108__I (.I(_01460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09109__A2 (.I(_01560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09110__A1 (.I(_01540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09115__S0 (.I(_01140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09115__S1 (.I(_01154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09116__A2 (.I(_01566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09117__A1 (.I(_01300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09118__B1 (.I(_01568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09119__A2 (.I(_01566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09120__A1 (.I(_01086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09121__A1 (.I(_01300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09122__A2 (.I(_01560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09123__A1 (.I(_01540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09128__S0 (.I(_01201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09128__S1 (.I(_01304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09129__S0 (.I(_01201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09129__S1 (.I(_01304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09130__A1 (.I(_01577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09131__A1 (.I(_01270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09132__I (.I(_01082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09136__I (.I(_01584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09137__I (.I(_01585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09138__A1 (.I(_01270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09138__A3 (.I(_01542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09139__A1 (.I(_01581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09140__I (.I(_01588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09141__A1 (.I(_01043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09141__A2 (.I(_01588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09142__I (.I(_01590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09145__B1 (.I(_01592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09150__S0 (.I(_01140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09150__S1 (.I(_01154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09152__A2 (.I(_01592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09152__B1 (.I(_01598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09157__I (.I(_01201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09158__I (.I(_01604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09159__I (.I(_01304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09160__I (.I(_01606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09161__S0 (.I(_01605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09161__S1 (.I(_01607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09162__A2 (.I(_01592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09164__I (.I(_01590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09165__I (.I(_01610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09169__S0 (.I(_01141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09169__S1 (.I(_01155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09170__B1 (.I(_01615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09175__S0 (.I(_01605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09175__S1 (.I(_01607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09181__S0 (.I(_01605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09181__S1 (.I(_01607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09182__I (.I(_01588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09183__I (.I(_01626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09189__S0 (.I(_01141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09189__S1 (.I(_01155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09190__B1 (.I(_01632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09192__I (.I(_01610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09196__S0 (.I(_01605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09196__S1 (.I(_01607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09202__I (.I(_01604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09203__I (.I(_01606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09204__S0 (.I(_01643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09204__S1 (.I(_01644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09210__S0 (.I(_01643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09210__S1 (.I(_01644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09211__I (.I(_01626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09217__I (.I(_01155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09218__S0 (.I(_01142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09218__S1 (.I(_01656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09219__B1 (.I(_01657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09221__I (.I(_01610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09225__S0 (.I(_01643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09225__S1 (.I(_01644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09226__A2 (.I(_01659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09231__S0 (.I(_01305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09231__S1 (.I(_01656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09232__A2 (.I(_01659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09232__B1 (.I(_01668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09237__S0 (.I(_01643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09237__S1 (.I(_01644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09238__I (.I(_01626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09239__A2 (.I(_01659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09244__I (.I(_01604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09245__I (.I(_01606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09246__S0 (.I(_01679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09246__S1 (.I(_01680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09247__A2 (.I(_01659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09249__I (.I(_01610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09253__I (.I(_01656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09255__S0 (.I(_01144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09255__S1 (.I(_01688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09256__A2 (.I(_01683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09256__B1 (.I(_01689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09261__S0 (.I(_01679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09261__S1 (.I(_01680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09262__A2 (.I(_01683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09266__S0 (.I(_01679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09266__S1 (.I(_01680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09267__I (.I(_01626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09268__A2 (.I(_01683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09268__B2 (.I(_01699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09270__A1 (.I(_01577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09270__B1 (.I(_01592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09275__I3 (.I(_01704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09275__S0 (.I(_01144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09276__A2 (.I(_01683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09276__B1 (.I(_01705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09276__B2 (.I(_01699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09281__I3 (.I(_01709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09281__S0 (.I(_01679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09281__S1 (.I(_01680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09282__B1 (.I(_01710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09282__B2 (.I(_01699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09287__S0 (.I(_01145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09287__S1 (.I(_01328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09288__B1 (.I(_01715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09288__B2 (.I(_01699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09293__S0 (.I(_01604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09293__S1 (.I(_01606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09295__A1 (.I(_01282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09296__I (.I(_01721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09298__I (.I(_01032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09299__A1 (.I(_01724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09299__A2 (.I(_01721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09303__A1 (.I(_01598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09305__A1 (.I(_01615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09306__I (.I(_01721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09307__I (.I(_01728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09309__I (.I(_01730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09312__A1 (.I(_01632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09314__I (.I(_01728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09315__I (.I(_01730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09318__A1 (.I(_01657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09320__I (.I(_01728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09321__I (.I(_01730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09322__A1 (.I(_01668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09322__A2 (.I(_01734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09322__B1 (.I(_01735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09323__A2 (.I(_01734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09323__B1 (.I(_01735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09324__A2 (.I(_01734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09324__B1 (.I(_01735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09325__A1 (.I(_01689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09325__A2 (.I(_01734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09325__B1 (.I(_01735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09326__I (.I(_01728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09327__I (.I(_01730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09330__A1 (.I(_01577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09331__A1 (.I(_01705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09332__A1 (.I(_01710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09333__A1 (.I(_01715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09336__I (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09338__I (.I(_01740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09339__I (.I(_01741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09340__I (.I(_01013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09341__I (.I(\filters.filt_1 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09346__I (.I(_01013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09347__I (.I(_01062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09348__I (.I(_01750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09349__I (.I(_01751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09350__I (.I(_01752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09351__A1 (.I(_01748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09351__B (.I(_01753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09352__A1 (.I(_01742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09353__I (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09354__I (.I(_01755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09355__I (.I(_01756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09356__I (.I(\filters.filt_2 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09361__I (.I(_01752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09362__A1 (.I(_01762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09363__A1 (.I(_01757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09364__I (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09366__I (.I(_01766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09367__I (.I(\filters.filt_3 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09373__A1 (.I(_01773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09374__A1 (.I(_01767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09375__I (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09377__I (.I(_01776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09378__A1 (.I(\filters.res_filt[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09379__A1 (.I(_01777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09380__I (.I(_01003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09381__I (.I(_01779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09382__I (.I(_01780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09383__I (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09384__A2 (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09385__I (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09386__A1 (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09387__I (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09388__I (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09393__A1 (.I(_01781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09397__A1 (.I(_01742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09398__I (.I(_01752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09400__A1 (.I(_01757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09402__A1 (.I(_01767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09403__A1 (.I(\filters.mode_vol[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09404__A1 (.I(_01777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09405__I (.I(_01017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09406__I (.I(_01800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09409__A1 (.I(\filters.lp ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09410__A1 (.I(_01801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09411__I (.I(_01006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09413__I (.I(_01806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09414__I (.I(_01751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09416__A1 (.I(\filters.bp ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09416__B (.I(_01809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09417__A1 (.I(_01807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09418__I (.I(net14));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09420__I (.I(_01812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09421__I (.I(_01813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09422__A1 (.I(\filters.hp ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09422__B (.I(_01809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09423__A1 (.I(_01814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09424__I (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09426__I (.I(_01817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09427__I (.I(_01818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09428__A1 (.I(\filters.mode_vol[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09428__B (.I(_01809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09429__A1 (.I(_01819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09430__I (.I(_01102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09431__I (.I(_01821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09432__I (.I(_01822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09440__A1 (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09440__A2 (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09443__I (.I(_01833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09444__A1 (.I(\channels.ctrl_reg2[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09444__A2 (.I(_01830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09448__A2 (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09452__A1 (.I(\channels.atk_dec2[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09452__B1 (.I(_01842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09452__B2 (.I(\channels.pw3[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09454__A1 (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09454__A2 (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09455__A2 (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09459__A1 (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09461__A1 (.I(\filters.cutoff_lut[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09461__B2 (.I(\filters.cutoff_lut[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09465__A2 (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09467__A1 (.I(\channels.freq1[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09467__B2 (.I(\channels.ctrl_reg1[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09469__A1 (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09470__A2 (.I(_01860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09472__A1 (.I(\channels.sus_rel3[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09472__B1 (.I(_01862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09472__B2 (.I(\channels.pw2[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09473__A1 (.I(_01852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09474__A1 (.I(_01748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09474__A2 (.I(_01844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09474__B2 (.I(\channels.pw2[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09476__I (.I(_01866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09479__A2 (.I(_01860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09481__B2 (.I(\channels.sus_rel2[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09481__C1 (.I(_01871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09481__C2 (.I(\channels.freq3[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09482__A3 (.I(_01865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09484__I (.I(_01874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09487__A1 (.I(\channels.ch3_env[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09491__I (.I(_01881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09492__B2 (.I(\channels.ctrl_reg3[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09493__A2 (.I(_01860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09497__A1 (.I(\channels.pw1[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09497__B2 (.I(\channels.freq1[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09503__A1 (.I(\channels.pw1[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09503__A2 (.I(_01891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09503__B2 (.I(\channels.freq2[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09506__B2 (.I(\channels.pw3[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09507__A2 (.I(_01860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09511__A2 (.I(_01899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09511__B2 (.I(\channels.atk_dec1[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09515__A1 (.I(\channels.sample3[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09515__A2 (.I(_01904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09515__B1 (.I(_01905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09515__B2 (.I(\clk_trg[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09516__A4 (.I(_01906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09517__I (.I(_01874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09519__A1 (.I(_01873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09519__A2 (.I(_01889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09519__B1 (.I(net22));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09520__A1 (.I(_01823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09521__A1 (.I(\channels.ctrl_reg2[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09521__A2 (.I(_01830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09522__A1 (.I(\channels.atk_dec2[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09522__B1 (.I(_01842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09522__B2 (.I(\channels.pw3[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09523__A1 (.I(\filters.cutoff_lut[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09523__B2 (.I(\filters.cutoff_lut[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09524__A1 (.I(\channels.freq1[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09524__B2 (.I(\channels.ctrl_reg1[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09525__A1 (.I(\channels.sus_rel3[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09525__B2 (.I(\channels.pw2[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09526__A1 (.I(_01913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09527__A1 (.I(_01762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09527__A2 (.I(_01844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09527__B2 (.I(\channels.pw2[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09528__B2 (.I(\channels.sus_rel2[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09528__C1 (.I(_01871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09528__C2 (.I(\channels.freq3[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09530__A1 (.I(\channels.ch3_env[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09531__B2 (.I(\channels.ctrl_reg3[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09532__A1 (.I(\channels.pw1[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09532__B2 (.I(\channels.freq1[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09534__A1 (.I(\channels.pw1[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09534__A2 (.I(_01891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09534__B2 (.I(\channels.freq2[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09535__B2 (.I(\channels.pw3[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09536__A2 (.I(_01899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09536__B2 (.I(\channels.atk_dec1[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09538__A1 (.I(_01927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09538__A2 (.I(_01904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09538__B1 (.I(_01905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09538__B2 (.I(\clk_trg[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09539__A4 (.I(_01928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09540__A1 (.I(_01919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09540__A2 (.I(_01923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09540__B1 (.I(net23));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09541__A1 (.I(_01823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09544__I (.I(_01932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09545__I (.I(_01874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09546__A1 (.I(\channels.ctrl_reg3[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09546__B1 (.I(_01862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09546__B2 (.I(\channels.pw2[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09549__A1 (.I(\channels.sus_rel2[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09549__B1 (.I(_01937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09549__B2 (.I(\channels.freq3[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09550__I (.I(_01904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09551__A1 (.I(_01773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09553__A1 (.I(\channels.pw1[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09553__B1 (.I(_01941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09553__B2 (.I(\channels.ctrl_reg1[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09555__A1 (.I(\filters.cutoff_lut[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09555__B1 (.I(_01943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09555__B2 (.I(\channels.sus_rel3[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09557__A1 (.I(\channels.sus_rel1[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09557__A2 (.I(_01899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09557__B1 (.I(_01939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09557__B2 (.I(\channels.sample3[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09560__A1 (.I(\channels.atk_dec1[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09561__A1 (.I(\channels.pw1[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09561__B2 (.I(\channels.freq2[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09562__A1 (.I(\channels.ctrl_reg2[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09562__B2 (.I(\channels.freq2[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09564__A1 (.I(\channels.pw3[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09564__A2 (.I(_01842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09564__B2 (.I(\channels.pw2[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09566__A1 (.I(\channels.ch3_env[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09566__B2 (.I(\channels.freq1[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09568__A1 (.I(\filters.cutoff_lut[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09568__A2 (.I(_01956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09568__B1 (.I(_01866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09568__B2 (.I(\channels.atk_dec3[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09569__A1 (.I(\channels.atk_dec2[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09569__B2 (.I(\channels.pw3[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09571__A1 (.I(\channels.freq1[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09571__A2 (.I(_01954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09571__B2 (.I(\channels.freq3[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09574__A1 (.I(_01933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09575__I (.I(_01943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09577__A1 (.I(\channels.sus_rel3[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09577__B1 (.I(_01964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09577__B2 (.I(\channels.sus_rel1[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09579__A1 (.I(\filters.res_filt[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09579__A2 (.I(_01844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09579__B2 (.I(\channels.freq2[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09580__A1 (.I(\filters.mode_vol[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09580__B2 (.I(\channels.sus_rel2[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09581__A1 (.I(\channels.ch3_env[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09581__B2 (.I(\channels.pw1[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09583__A1 (.I(\channels.pw3[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09583__B1 (.I(_01970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09583__B2 (.I(\channels.freq1[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09585__A1 (.I(\channels.atk_dec2[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09587__A1 (.I(\channels.pw1[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09587__A2 (.I(_01891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09588__A1 (.I(\channels.freq3[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09590__A1 (.I(\channels.ctrl_reg1[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09590__A2 (.I(_01941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09590__B2 (.I(_01977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09591__A1 (.I(_01874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09592__A1 (.I(\channels.ctrl_reg2[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09592__B2 (.I(\channels.ctrl_reg3[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09593__A1 (.I(\channels.pw2[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09593__B2 (.I(\channels.atk_dec1[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09594__A1 (.I(\channels.atk_dec3[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09594__B2 (.I(\channels.pw3[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09595__A1 (.I(\filters.cutoff_lut[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09595__A2 (.I(_01956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09595__B1 (.I(_01954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09595__B2 (.I(\channels.freq1[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09597__B1 (.I(_01862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09597__B2 (.I(\channels.pw2[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09599__A2 (.I(net25));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09600__A1 (.I(_01933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09601__I (.I(_01956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09602__A1 (.I(\filters.cutoff_lut[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09603__A1 (.I(\channels.sus_rel3[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09603__B2 (.I(\channels.freq1[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09604__I (.I(_01866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09605__I (.I(_01833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09607__A2 (.I(_01989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09608__A1 (.I(\channels.ctrl_reg2[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09608__B2 (.I(\channels.atk_dec2[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09611__A1 (.I(\channels.pw2[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09611__B2 (.I(\channels.freq2[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09612__I (.I(_01881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09613__A1 (.I(\channels.freq3[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09613__A2 (.I(_01937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09613__B2 (.I(\channels.ctrl_reg3[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09615__A1 (.I(\channels.sus_rel2[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09617__I (.I(_01941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09618__A1 (.I(\channels.pw1[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09618__B2 (.I(\channels.ctrl_reg1[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09620__I (.I(_01844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09621__B1 (.I(_01939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09621__B2 (.I(\channels.sample3[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09623__A1 (.I(\channels.ch3_env[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09623__B2 (.I(\channels.atk_dec1[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09624__I (.I(_01954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09626__A1 (.I(\channels.freq1[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09626__B2 (.I(\channels.pw3[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09628__A1 (.I(\filters.lp ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09628__B1 (.I(_01964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09628__B2 (.I(\channels.sus_rel1[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09629__A1 (.I(_02008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09631__A2 (.I(net26));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09631__B (.I(_01809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09632__A2 (.I(_02017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09633__A1 (.I(\filters.cutoff_lut[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09634__A1 (.I(\channels.sus_rel3[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09634__B1 (.I(_01970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09634__B2 (.I(\channels.freq1[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09636__A2 (.I(_02019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09637__A1 (.I(\channels.ctrl_reg2[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09637__B2 (.I(\channels.atk_dec2[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09638__A1 (.I(\channels.pw2[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09638__B2 (.I(\channels.freq2[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09639__A2 (.I(_01937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09639__B2 (.I(\channels.ctrl_reg3[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09640__A1 (.I(\channels.sus_rel2[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09641__A1 (.I(\channels.pw1[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09641__B2 (.I(\channels.ctrl_reg1[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09644__A1 (.I(\filters.res_filt[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09644__B1 (.I(_01939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09644__B2 (.I(_02029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09645__A1 (.I(\channels.ch3_env[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09645__B2 (.I(\channels.atk_dec1[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09646__A1 (.I(\channels.freq1[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09646__B2 (.I(\channels.pw3[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09647__A1 (.I(\filters.bp ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09647__B1 (.I(_01964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09647__B2 (.I(\channels.sus_rel1[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09648__A1 (.I(_02030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09651__A2 (.I(net27));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09651__B (.I(_02036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09652__A2 (.I(_02035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09653__A1 (.I(\filters.cutoff_lut[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09654__A1 (.I(\channels.sus_rel3[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09654__A2 (.I(_01943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09654__B1 (.I(_01970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09654__B2 (.I(\channels.freq1[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09656__A2 (.I(_02038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09657__A1 (.I(\channels.ctrl_reg2[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09657__B2 (.I(\channels.atk_dec2[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09658__B2 (.I(\channels.freq2[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09659__A2 (.I(_01871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09659__B2 (.I(\channels.ctrl_reg3[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09660__A1 (.I(\channels.sus_rel2[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09661__A1 (.I(\channels.pw1[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09661__B2 (.I(\channels.ctrl_reg1[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09663__A1 (.I(\filters.res_filt[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09663__B1 (.I(_01939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09663__B2 (.I(\channels.sample3[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09664__A1 (.I(\channels.ch3_env[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09664__B2 (.I(\channels.atk_dec1[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09665__A1 (.I(\channels.freq1[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09665__B2 (.I(\channels.pw3[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09666__A1 (.I(\filters.hp ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09666__B1 (.I(_01899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09666__B2 (.I(\channels.sus_rel1[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09667__A1 (.I(_02048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09669__A2 (.I(net28));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09669__B (.I(_02036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09670__A2 (.I(_02053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09672__I (.I(\channels.sample3[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09673__A1 (.I(\channels.ctrl_reg2[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09673__A2 (.I(_01830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09673__B1 (.I(_01904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09673__B2 (.I(_02056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09674__A1 (.I(\channels.atk_dec1[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09674__B (.I(_01905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09676__A1 (.I(\channels.sus_rel3[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09676__B1 (.I(_01964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09676__B2 (.I(\channels.sus_rel1[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09677__A1 (.I(\channels.freq1[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09677__B2 (.I(\channels.sus_rel2[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09678__A1 (.I(\filters.mode_vol[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09679__A1 (.I(\channels.freq2[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09679__B2 (.I(\channels.freq1[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09680__A1 (.I(\channels.atk_dec2[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09680__B1 (.I(_01937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09680__B2 (.I(\channels.freq3[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09682__A1 (.I(\channels.ctrl_reg3[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09682__B2 (.I(\channels.ctrl_reg1[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09683__A1 (.I(\filters.cutoff_lut[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09683__B2 (.I(\channels.ch3_env[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09684__A1 (.I(\filters.res_filt[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09685__A1 (.I(\channels.pw1[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09688__A1 (.I(net29));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09688__B (.I(_02036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09689__A2 (.I(_02071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09690__A1 (.I(_01781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09690__A2 (.I(_01970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09693__A1 (.I(\channels.freq1[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09693__B (.I(_02036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09694__A1 (.I(_01742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09696__A1 (.I(\channels.freq1[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09697__A1 (.I(_01757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09698__A1 (.I(\channels.freq1[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09699__A1 (.I(_01767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09700__A1 (.I(\channels.freq1[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09701__A1 (.I(_01777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09704__A1 (.I(\channels.freq1[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09705__A1 (.I(_01801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09707__A1 (.I(\channels.freq1[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09708__A1 (.I(_01807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09709__A1 (.I(\channels.freq1[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09710__A1 (.I(_01814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09711__A1 (.I(\channels.freq1[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09712__A1 (.I(_01819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09713__I (.I(_01780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09714__A1 (.I(_02088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09714__A2 (.I(_01891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09717__A1 (.I(\channels.pw1[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09718__A1 (.I(_01742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09719__I (.I(_01751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09721__A1 (.I(\channels.pw1[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09722__A1 (.I(_01757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09723__A1 (.I(\channels.pw1[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09724__A1 (.I(_01767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09725__I (.I(\channels.pw1[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09726__I (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09727__A1 (.I(_02098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09728__I (.I(_01062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09730__I (.I(_02101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09732__C (.I(_02103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09734__I (.I(_02104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09735__A1 (.I(_01781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09735__A2 (.I(_01941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09736__I (.I(_02106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09737__I (.I(_02106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09738__A1 (.I(\channels.ctrl_reg1[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09740__I (.I(_01756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09741__A1 (.I(\channels.ctrl_reg1[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09742__A1 (.I(_02110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09743__I (.I(_01766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09745__A1 (.I(\channels.ctrl_reg1[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09745__B (.I(_02113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09746__A1 (.I(_02112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09747__A1 (.I(\channels.ctrl_reg1[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09747__B (.I(_02113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09748__A1 (.I(_01777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09749__I (.I(_02106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09750__I (.I(_02106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09751__A1 (.I(\channels.ctrl_reg1[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09751__B (.I(_02113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09752__A1 (.I(_01801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09753__A1 (.I(\channels.ctrl_reg1[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09753__B (.I(_02113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09754__A1 (.I(_01807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09756__A1 (.I(\channels.ctrl_reg1[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09756__B (.I(_02120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09757__A1 (.I(_01814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09758__A1 (.I(\channels.ctrl_reg1[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09758__B (.I(_02120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09759__A1 (.I(_01819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09760__I (.I(_01780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09764__A1 (.I(\channels.atk_dec1[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09764__B (.I(_02120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09766__A1 (.I(\channels.atk_dec1[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09766__B (.I(_02120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09767__A1 (.I(_02110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09769__A1 (.I(\channels.atk_dec1[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09770__A1 (.I(_02112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09771__I (.I(_01776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09772__A1 (.I(\channels.atk_dec1[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09773__A1 (.I(_02131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09776__A1 (.I(\channels.atk_dec1[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09777__A1 (.I(_01801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09778__A1 (.I(\channels.atk_dec1[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09779__A1 (.I(_01807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09780__I (.I(_01751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09782__A1 (.I(\channels.atk_dec1[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09783__A1 (.I(_01814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09784__A1 (.I(\channels.atk_dec1[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09785__A1 (.I(_01819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09792__A1 (.I(_02110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09794__A1 (.I(\channels.sus_rel1[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09795__A1 (.I(_02112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09796__A1 (.I(\channels.sus_rel1[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09797__A1 (.I(_02131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09798__I (.I(_01017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09799__I (.I(_02149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09802__A1 (.I(\channels.sus_rel1[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09803__A1 (.I(_02150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09805__I (.I(_02154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09806__A1 (.I(\channels.sus_rel1[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09807__A1 (.I(_02155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09808__I (.I(_01813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09810__A1 (.I(\channels.sus_rel1[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09812__I (.I(_01818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09813__A1 (.I(\channels.sus_rel1[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09814__A1 (.I(_02160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09818__A1 (.I(\channels.freq2[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09820__A1 (.I(\channels.freq2[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09821__A1 (.I(_02110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09823__A1 (.I(\channels.freq2[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09824__A1 (.I(_02112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09825__A1 (.I(\channels.freq2[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09826__A1 (.I(_02131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09829__A1 (.I(\channels.freq2[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09830__A1 (.I(_02150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09831__A1 (.I(\channels.freq2[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09832__A1 (.I(_02155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09833__I (.I(_01750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09834__I (.I(_02174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09836__A1 (.I(\channels.freq2[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09838__A1 (.I(\channels.freq2[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09839__A1 (.I(_02160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09840__I (.I(_02104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09841__A1 (.I(_02088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09841__A2 (.I(_01862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09844__A1 (.I(\channels.pw2[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09845__A1 (.I(_02179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09846__I (.I(_01755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09847__I (.I(_02184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09848__A1 (.I(\channels.pw2[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09851__I (.I(_02187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09853__A1 (.I(\channels.pw2[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09855__I (.I(\channels.pw2[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09856__A1 (.I(_02098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09857__C (.I(_02103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09858__A2 (.I(_01830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09861__A1 (.I(\channels.ctrl_reg2[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09862__A1 (.I(_02179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09863__A1 (.I(\channels.ctrl_reg2[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09865__A1 (.I(\channels.ctrl_reg2[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09868__A1 (.I(\channels.ctrl_reg2[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09869__A1 (.I(_02131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09872__A1 (.I(\channels.ctrl_reg2[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09873__A1 (.I(_02150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09874__A1 (.I(\channels.ctrl_reg2[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09875__A1 (.I(_02155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09876__A1 (.I(\channels.ctrl_reg2[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09879__A1 (.I(\channels.ctrl_reg2[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09880__A1 (.I(_02160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09881__I (.I(_01779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09883__I (.I(_02209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09884__I (.I(_02209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09885__A1 (.I(\channels.atk_dec2[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09886__A1 (.I(_02179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09887__A1 (.I(\channels.atk_dec2[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09889__A1 (.I(\channels.atk_dec2[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09891__I (.I(_01776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09892__I (.I(_02174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09894__A1 (.I(\channels.atk_dec2[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09895__A1 (.I(_02215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09896__I (.I(_02209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09897__I (.I(_02209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09898__A1 (.I(\channels.atk_dec2[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09899__A1 (.I(_02150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09900__A1 (.I(\channels.atk_dec2[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09901__A1 (.I(_02155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09902__A1 (.I(\channels.atk_dec2[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09905__A1 (.I(\channels.atk_dec2[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09906__A1 (.I(_02160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09908__I (.I(_02226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09909__I (.I(_02226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09910__A1 (.I(\channels.sus_rel2[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09911__A1 (.I(_02179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09912__A1 (.I(\channels.sus_rel2[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09914__A1 (.I(\channels.sus_rel2[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09917__A1 (.I(\channels.sus_rel2[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09917__B (.I(_02232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09918__A1 (.I(_02215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09919__I (.I(_02149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09920__I (.I(_02226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09921__I (.I(_02226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09922__A1 (.I(\channels.sus_rel2[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09922__B (.I(_02232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09923__A1 (.I(_02234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09924__I (.I(_02154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09925__A1 (.I(\channels.sus_rel2[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09925__B (.I(_02232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09926__A1 (.I(_02238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09927__I (.I(_01813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09928__A1 (.I(\channels.sus_rel2[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09928__B (.I(_02232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09929__A1 (.I(_02240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09930__I (.I(_01818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09932__A1 (.I(\channels.sus_rel2[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09932__B (.I(_02243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09933__A1 (.I(_02242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09934__I (.I(_02104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09935__A2 (.I(_01833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09938__B (.I(_02243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09939__A1 (.I(_02245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09940__I (.I(_02184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09941__B (.I(_02243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09942__A1 (.I(_02250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09943__I (.I(_02187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09944__A1 (.I(\channels.freq3[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09944__B (.I(_02243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09945__A1 (.I(_02252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09946__I (.I(_02174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09947__I (.I(_02254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09949__A1 (.I(_02215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09953__A1 (.I(_02234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09955__A1 (.I(_02238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09957__A1 (.I(_02240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09958__I (.I(_02254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09960__A1 (.I(_02242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09961__A1 (.I(_01781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09961__A2 (.I(_01842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09964__A1 (.I(\channels.pw3[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09964__A2 (.I(_02266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09965__A1 (.I(_02245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09965__A2 (.I(_02265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09966__A1 (.I(\channels.pw3[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09966__A2 (.I(_02266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09967__A1 (.I(_02250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09967__A2 (.I(_02265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09968__A1 (.I(\channels.pw3[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09968__A2 (.I(_02266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09969__A1 (.I(_02252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09969__A2 (.I(_02265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09970__I (.I(\channels.pw3[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09971__A1 (.I(_02098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09971__A2 (.I(_02266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09972__I (.I(_02101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09973__I (.I(_02272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09974__A2 (.I(_02265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09974__C (.I(_02273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09975__A2 (.I(_01881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09978__I (.I(_02254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09979__A1 (.I(\channels.ctrl_reg3[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09980__A1 (.I(_02245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09981__A1 (.I(\channels.ctrl_reg3[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09982__A1 (.I(_02250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09983__A1 (.I(\channels.ctrl_reg3[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09984__A1 (.I(_02252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09985__A1 (.I(\channels.ctrl_reg3[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09986__A1 (.I(_02215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09989__I (.I(_02254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09990__A1 (.I(\channels.ctrl_reg3[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09991__A1 (.I(_02234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09992__A1 (.I(\channels.ctrl_reg3[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09993__A1 (.I(_02238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09994__A1 (.I(\channels.ctrl_reg3[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09995__A1 (.I(_02240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09996__A1 (.I(\channels.ctrl_reg3[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09997__A1 (.I(_02242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09998__I (.I(_01779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09999__A1 (.I(_02289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10000__I (.I(_02290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10001__I (.I(_02290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10002__I (.I(_02174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10003__I (.I(_02293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10005__A1 (.I(_02245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10007__A1 (.I(_02250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10008__A1 (.I(\channels.atk_dec3[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10009__A1 (.I(_02252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10012__A1 (.I(\channels.atk_dec3[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10013__A1 (.I(_02299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10014__I (.I(_02290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10015__I (.I(_02290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10016__I (.I(_02293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10018__A1 (.I(_02234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10020__A1 (.I(_02238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10022__A1 (.I(_02240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10024__A1 (.I(_02242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10025__I (.I(_02104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10026__A1 (.I(_02289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10026__A2 (.I(_01943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10029__I (.I(_02293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10030__A1 (.I(\channels.sus_rel3[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10031__A1 (.I(_02308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10032__I (.I(_02184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10033__A1 (.I(\channels.sus_rel3[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10034__A1 (.I(_02314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10035__I (.I(_02187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10036__A1 (.I(\channels.sus_rel3[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10037__A1 (.I(_02316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10038__A1 (.I(\channels.sus_rel3[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10039__A1 (.I(_02299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10040__I (.I(_02149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10043__I (.I(_02293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10044__A1 (.I(\channels.sus_rel3[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10045__A1 (.I(_02319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10046__I (.I(_02154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10047__A1 (.I(\channels.sus_rel3[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10048__A1 (.I(_02324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10049__I (.I(_01813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10050__A1 (.I(\channels.sus_rel3[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10051__A1 (.I(_02326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10052__I (.I(_01818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10053__A1 (.I(\channels.sus_rel3[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10054__A1 (.I(_02328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10055__A1 (.I(_02289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10055__A2 (.I(_01956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10056__I (.I(_02330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10057__I (.I(_02330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10058__I (.I(_01750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10060__I (.I(_02334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10061__A1 (.I(\filters.cutoff_lut[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10062__A1 (.I(_02308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10063__A1 (.I(\filters.cutoff_lut[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10064__A1 (.I(_02314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10065__A1 (.I(\filters.cutoff_lut[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10066__A1 (.I(_02316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10067__A1 (.I(\filters.cutoff_lut[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10068__A1 (.I(_02299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10069__I (.I(_02330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10070__I (.I(_02330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10071__I (.I(_02334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10072__A1 (.I(\filters.cutoff_lut[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10073__A1 (.I(_02319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10074__A1 (.I(\filters.cutoff_lut[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10075__A1 (.I(_02324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10076__A1 (.I(\filters.cutoff_lut[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10077__A1 (.I(_02326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10078__A1 (.I(\filters.cutoff_lut[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10079__A1 (.I(_02328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10083__A1 (.I(_01933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10084__I (.I(\clk_trg[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10085__A1 (.I(_02088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10085__A2 (.I(_01905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10086__A1 (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10086__A2 (.I(_02351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10087__I (.I(_01724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10089__A2 (.I(_02351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10089__C (.I(_02354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10090__A1 (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10090__A2 (.I(_02351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10091__A2 (.I(_02351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10091__C (.I(_02354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10092__I (.I(_01082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10093__A1 (.I(_01070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10093__A2 (.I(_02356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10096__I (.I(_01085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10098__A2 (.I(_01245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10099__A1 (.I(_02359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10100__I (.I(_01282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10101__A1 (.I(_01070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10101__A2 (.I(_02363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10102__I (.I(_02364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10103__I (.I(_02365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10104__A2 (.I(_01230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10105__A1 (.I(_02366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10106__A2 (.I(_01560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10107__A1 (.I(_01540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10108__A2 (.I(\channels.ctrl_reg2[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10109__A2 (.I(\channels.ctrl_reg3[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10109__B1 (.I(\channels.ctrl_reg1[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10111__I (.I(_02371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10112__A1 (.I(\channels.ctrl_reg2[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10112__A2 (.I(\channels.ring_outs[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10113__A1 (.I(\channels.ctrl_reg3[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10113__A2 (.I(\channels.ring_outs[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10114__A1 (.I(\channels.ctrl_reg1[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10114__A2 (.I(\channels.ring_outs[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10116__A2 (.I(_02376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10117__I (.I(_02377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10118__A1 (.I(_01527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10119__A1 (.I(\channels.ctrl_reg1[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10119__A2 (.I(_01286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10120__A1 (.I(\channels.ctrl_reg3[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10120__B2 (.I(\channels.ctrl_reg2[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10121__I (.I(_02381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10122__A1 (.I(\channels.ctrl_reg3[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10123__A1 (.I(\channels.ctrl_reg2[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10123__B1 (.I(_01286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10123__B2 (.I(\channels.ctrl_reg1[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10125__I (.I(_02385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10126__A1 (.I(_01632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10127__A1 (.I(_01534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10130__A3 (.I(\channels.pw3[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10131__A2 (.I(\channels.pw2[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10132__A1 (.I(\channels.pw1[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10137__A3 (.I(\channels.pw2[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10138__A3 (.I(\channels.pw3[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10139__A1 (.I(\channels.pw1[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10141__S0 (.I(_01495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10141__S1 (.I(_01496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10142__A1 (.I(_01085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10142__B2 (.I(_02402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10143__I (.I(_01555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10145__A3 (.I(\channels.pw3[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10146__A2 (.I(\channels.pw2[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10147__A1 (.I(\channels.pw1[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10149__A3 (.I(\channels.pw2[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10150__A3 (.I(\channels.pw3[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10151__A1 (.I(\channels.pw1[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10155__A1 (.I(_01566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10160__A1 (.I(_01555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10160__B2 (.I(_01550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10170__A1 (.I(\channels.pw1[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10171__A1 (.I(_01541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10173__I (.I(\channels.pw1[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10175__A3 (.I(\channels.pw3[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10176__A2 (.I(\channels.pw2[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10177__C (.I(_01527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10178__I (.I(\channels.pw1[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10179__A3 (.I(\channels.pw3[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10180__A2 (.I(\channels.pw2[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10181__A2 (.I(_01286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10181__C (.I(_01520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10184__A3 (.I(\channels.pw3[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10185__A1 (.I(\channels.pw1[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10186__A1 (.I(_01533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10187__A3 (.I(\channels.pw2[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10188__A1 (.I(\channels.pw1[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10189__A1 (.I(_01527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10192__A1 (.I(_01541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10192__C2 (.I(_01533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10193__I (.I(\channels.pw2[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10195__A2 (.I(_02455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10195__A3 (.I(\channels.pw3[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10196__A1 (.I(\channels.pw1[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10197__A2 (.I(_01099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10199__A3 (.I(\channels.pw2[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10200__A2 (.I(_02455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10200__A3 (.I(\channels.pw3[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10201__A1 (.I(\channels.pw1[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10202__A1 (.I(_01469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10203__A3 (.I(\channels.pw3[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10204__A2 (.I(\channels.pw1[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10205__A2 (.I(\channels.pw2[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10206__A1 (.I(_01481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10207__B (.I(_01481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10209__I (.I(\channels.pw2[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10210__A2 (.I(_02455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10210__A3 (.I(\channels.pw3[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10211__A1 (.I(\channels.pw1[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10212__A2 (.I(_01099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10213__A2 (.I(_02473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10215__A1 (.I(_01541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10215__B2 (.I(_01533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10217__A3 (.I(\channels.pw2[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10218__A1 (.I(\channels.pw1[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10219__A1 (.I(_01520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10220__A2 (.I(_02473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10227__A1 (.I(_01481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10229__A1 (.I(_01510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10229__A2 (.I(_02473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10231__B (.I(_01469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10234__A2 (.I(\channels.ctrl_reg2[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10236__A2 (.I(\channels.ctrl_reg3[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10236__B1 (.I(\channels.ctrl_reg1[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10238__A1 (.I(_02484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10238__A2 (.I(_02498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10240__I (.I(_02500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10242__I2 (.I(\channels.ch3_env[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10242__S0 (.I(_01145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10242__S1 (.I(_01159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10243__I (.I(_02503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10245__A1 (.I(_02502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10245__A2 (.I(_02505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10246__A1 (.I(_02484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10246__A2 (.I(_02498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10247__I (.I(_02507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10249__A1 (.I(_01497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10250__A1 (.I(_01508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10250__A2 (.I(_02381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10252__I (.I(_02512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10254__I (.I(\channels.ch3_env[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10257__I (.I(_01141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10261__A1 (.I(_01688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10262__A3 (.I(_02522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10264__A1 (.I(_01482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10265__A1 (.I(_01497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10267__I (.I(_02527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10268__I (.I(_01656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10269__I (.I(\channels.ch3_env[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10270__A1 (.I(_01305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10275__I (.I(_02535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10279__A1 (.I(_01470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10281__A1 (.I(_01482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10283__I2 (.I(\channels.ch3_env[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10284__A2 (.I(_02543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10284__A3 (.I(_02544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10288__A1 (.I(_01521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10288__A2 (.I(_02377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10289__I (.I(_02371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10290__A1 (.I(_01615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10290__A2 (.I(_02385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10291__A1 (.I(_01528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10292__A1 (.I(_02484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10292__A2 (.I(_02498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10293__I (.I(_02553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10295__I (.I(\channels.ch3_env[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10296__A1 (.I(_01307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10297__A1 (.I(_01307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10298__S (.I(_01144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10299__A1 (.I(_01328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10300__A1 (.I(_01328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10301__I (.I(_02561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10302__A1 (.I(_02555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10307__A1 (.I(_01470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10309__I (.I(\channels.ch3_env[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10312__S (.I(_01142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10315__I (.I(_02575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10316__A2 (.I(_02569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10317__I (.I(\channels.ch3_env[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10322__A1 (.I(_01688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10323__A2 (.I(_02543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10325__A1 (.I(_01510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10325__A2 (.I(_02377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10326__A1 (.I(_01598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10326__A2 (.I(_02385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10327__A1 (.I(_01521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10327__A2 (.I(_02381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10328__A1 (.I(_02484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10328__A2 (.I(_02498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10330__A1 (.I(_02522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10330__A2 (.I(_02590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10331__I (.I(_02507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10332__A2 (.I(_02535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10333__I (.I(_02544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10339__I (.I(_02569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10342__A3 (.I(_02602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10346__I (.I(_02503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10347__A1 (.I(_02502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10347__A2 (.I(_02607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10356__A2 (.I(_02502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10358__A1 (.I(_01534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10359__A1 (.I(_01657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10360__A1 (.I(_01542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10362__I (.I(_02622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10364__A2 (.I(_02624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10369__I (.I(_02543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10371__I (.I(\channels.ch3_env[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10372__A1 (.I(_01305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10378__A2 (.I(_02569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10378__A3 (.I(_02638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10380__I (.I(_02522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10382__A1 (.I(_02642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10382__A2 (.I(_02555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10384__I (.I(_02590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10392__A1 (.I(_02555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10392__A2 (.I(_02503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10393__A3 (.I(_02642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10396__I (.I(_02544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10397__A2 (.I(_02657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10397__A3 (.I(_02569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10401__I (.I(_02561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10402__A1 (.I(_02662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10414__A3 (.I(_02662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10416__A2 (.I(_02676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10419__A1 (.I(_02607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10426__I (.I(_02686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10427__A3 (.I(_02687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10436__A3 (.I(_02686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10437__A3 (.I(_02607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10442__I (.I(_02505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10444__A1 (.I(_01162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10445__A1 (.I(_01162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10447__A2 (.I(_02707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10448__A3 (.I(_02703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10449__I (.I(_02642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10450__I (.I(_02505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10451__A2 (.I(_02527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10453__B1 (.I(_02711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10454__A2 (.I(_02710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10459__A1 (.I(_01164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10460__A1 (.I(_01164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10461__A2 (.I(_02721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10462__A2 (.I(_02703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10476__A1 (.I(_02703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10476__A3 (.I(_02624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10487__A2 (.I(_02543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10487__A3 (.I(_02638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10489__A1 (.I(_02507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10489__A2 (.I(_02512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10490__A1 (.I(_01688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10492__A2 (.I(_02752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10501__A2 (.I(_02754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10505__A1 (.I(_02662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10508__A1 (.I(_01542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10511__A1 (.I(_01668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10512__A1 (.I(_01550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10517__A2 (.I(_02777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10523__I (.I(_01089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10524__A1 (.I(\channels.sample3[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10525__A1 (.I(_02359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10525__A2 (.I(_02783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10531__A1 (.I(_02686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10531__A2 (.I(_02624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10535__A2 (.I(_02754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10536__A2 (.I(_02754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10547__A2 (.I(_02590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10550__A1 (.I(_02522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10550__A2 (.I(_02622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10551__A1 (.I(_02544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10552__A1 (.I(_02535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10552__A2 (.I(_02500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10558__A1 (.I(_02561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10560__A1 (.I(_01550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10561__A1 (.I(_01689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10562__A1 (.I(_01556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10564__I (.I(_02823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10565__A1 (.I(_02607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10572__A1 (.I(\channels.sample3[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10573__A1 (.I(_02359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10573__A2 (.I(_02831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10579__A1 (.I(_02687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10579__A2 (.I(_02777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10580__I (.I(_02703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10582__A1 (.I(_02839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10582__A3 (.I(_02840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10589__B1 (.I(_02847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10590__A4 (.I(_02847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10594__A1 (.I(_02575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10601__A2 (.I(_02500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10602__A2 (.I(_02622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10608__A2 (.I(_02823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10610__A1 (.I(_01556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10611__A1 (.I(_01705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10612__A1 (.I(_02402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10614__I (.I(_02872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10622__A1 (.I(\channels.sample3[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10623__A1 (.I(_02359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10623__A2 (.I(_02880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10631__A1 (.I(_02687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10631__A2 (.I(_02840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10633__A1 (.I(_02839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10633__A3 (.I(_02890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10643__A1 (.I(_02590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10644__A1 (.I(_02553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10644__A2 (.I(_02575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10650__A1 (.I(_02642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10650__A2 (.I(_02823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10651__A1 (.I(_02657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10651__A2 (.I(_02622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10660__A1 (.I(_02662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10660__A2 (.I(_02872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10662__A1 (.I(_02402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10663__A1 (.I(_01715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10664__A1 (.I(_01085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10666__A1 (.I(_02505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10666__A2 (.I(_02923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10675__A1 (.I(\channels.sample3[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10676__A2 (.I(_02932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10682__I (.I(_02923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10684__A1 (.I(_02839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10684__A3 (.I(_02940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10691__A1 (.I(_02686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10691__A2 (.I(_02923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10696__A1 (.I(_02602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10697__A1 (.I(_02555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10697__A2 (.I(_02638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10703__A1 (.I(_02710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10704__I (.I(_02657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10705__A2 (.I(_02777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10706__A1 (.I(_02676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10718__I (.I(_02974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10719__A1 (.I(\channels.sample3[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10720__A2 (.I(_02973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10737__A1 (.I(_02602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10738__I (.I(_02638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10739__A1 (.I(_02502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10744__A1 (.I(_02710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10744__A2 (.I(_02923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10745__A1 (.I(_02657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10745__A2 (.I(_02823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10746__A1 (.I(_02676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10746__A2 (.I(_02872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10758__A1 (.I(_01927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10759__A2 (.I(_03013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10773__I (.I(_02602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10774__A2 (.I(_02840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10775__A1 (.I(_02624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10777__A2 (.I(_02777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10784__I (.I(_02676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10785__A1 (.I(_03039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10798__A1 (.I(\channels.sample3[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10799__A2 (.I(_03052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10810__A2 (.I(_02872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10827__A1 (.I(_01977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10828__A2 (.I(_03080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10836__A2 (.I(_02840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10837__A2 (.I(_02890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10844__A2 (.I(_02940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10852__I (.I(_02974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10853__A1 (.I(\channels.sample3[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10854__A2 (.I(_03104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10861__A2 (.I(_02890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10862__A2 (.I(_02940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10871__A1 (.I(_02029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10872__A2 (.I(_03122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10879__A1 (.I(_03128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10879__A2 (.I(_02890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10881__A1 (.I(_03131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10881__A2 (.I(_02940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10886__A1 (.I(\channels.sample3[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10887__A2 (.I(_03136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10892__A1 (.I(_02056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10893__A1 (.I(_03138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10893__A2 (.I(_03141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10894__I (.I(_01104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10895__A1 (.I(\channels.sample2[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10896__A1 (.I(_02366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10896__A2 (.I(_02783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10897__A1 (.I(\channels.sample2[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10898__A1 (.I(_02366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10898__A2 (.I(_02831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10899__A1 (.I(\channels.sample2[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10900__A1 (.I(_02366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10900__A2 (.I(_02880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10901__I (.I(_02365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10902__A1 (.I(\channels.sample2[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10903__A2 (.I(_02932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10905__I (.I(_03149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10906__A1 (.I(\channels.sample2[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10907__A2 (.I(_02973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10908__A1 (.I(\channels.sample2[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10909__A2 (.I(_03013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10910__A1 (.I(\channels.sample2[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10911__A2 (.I(_03052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10912__I (.I(_02365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10913__A1 (.I(\channels.sample2[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10914__A2 (.I(_03080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10915__I (.I(_03149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10916__A1 (.I(\channels.sample2[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10916__A2 (.I(_03156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10917__A2 (.I(_03104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10918__A1 (.I(\channels.sample2[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10918__A2 (.I(_03156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10919__A2 (.I(_03122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10920__A1 (.I(\channels.sample2[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10920__A2 (.I(_03156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10921__A2 (.I(_03136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10922__I (.I(_02365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10923__A1 (.I(\channels.sample2[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10923__A2 (.I(_03156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10924__A2 (.I(_03141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10925__I (.I(_01321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10926__A1 (.I(\channels.sample1[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10926__A2 (.I(_01560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10927__A2 (.I(_02783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10928__I (.I(_01460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10929__A1 (.I(\channels.sample1[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10930__A2 (.I(_02831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10931__A1 (.I(\channels.sample1[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10932__A2 (.I(_02880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10933__A1 (.I(\channels.sample1[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10934__A2 (.I(_02932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10935__I (.I(_01320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10936__A1 (.I(\channels.sample1[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10937__A2 (.I(_02973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10938__I (.I(_01460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10939__A1 (.I(\channels.sample1[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10940__A2 (.I(_03013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10941__A1 (.I(\channels.sample1[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10942__A2 (.I(_03052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10943__A1 (.I(\channels.sample1[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10944__A2 (.I(_03080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10945__I (.I(_01320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10946__A1 (.I(\channels.sample1[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10947__A2 (.I(_03104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10948__A1 (.I(\channels.sample1[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10948__A2 (.I(_01261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10949__A2 (.I(_03122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10950__A1 (.I(\channels.sample1[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10950__A2 (.I(_01261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10951__A2 (.I(_03136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10952__A1 (.I(\channels.sample1[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10952__A2 (.I(_01261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10953__A2 (.I(_03141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10960__I (.I(_03184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10961__I (.I(_03185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10963__I (.I(_03187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10974__A2 (.I(_03194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10975__I (.I(_03199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10980__A1 (.I(_03202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10980__A2 (.I(_03204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10981__A2 (.I(_03205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10982__I (.I(_03206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10983__B (.I(_03200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10984__A2 (.I(_03205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10989__I (.I(_03204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10991__I (.I(_03215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10997__I (.I(_03221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11002__A1 (.I(\filters.lp ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11002__A2 (.I(_03226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11012__A1 (.I(_03204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11012__A2 (.I(_03215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11015__A1 (.I(\filters.hp ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11015__A2 (.I(_03236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11015__B2 (.I(\filters.bp ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11015__C (.I(_03239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11016__A1 (.I(_01069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11021__A3 (.I(_03243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11021__B1 (.I(_03245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11028__B (.I(_03251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11033__A2 (.I(_03187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11033__B (.I(_03256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11033__C (.I(_03206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11034__A1 (.I(\filters.high[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11040__A1 (.I(_03243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11040__B1 (.I(_03245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11040__B2 (.I(_03263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11044__B (.I(_03263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11048__I (.I(_03270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11051__B (.I(_03273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11051__C (.I(_03206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11052__A1 (.I(\filters.high[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11063__B (.I(_03284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11067__B (.I(_03288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11067__C (.I(_03206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11068__A1 (.I(\filters.high[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11079__B (.I(_03299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11082__A1 (.I(\filters.low[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11082__B (.I(_03302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11095__B (.I(_03314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11097__I (.I(_03316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11098__A1 (.I(_03310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11098__B (.I(_03317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11099__A1 (.I(\filters.high[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11112__B (.I(_03330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11115__A1 (.I(_03329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11115__B (.I(_03333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11117__A1 (.I(\filters.high[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11119__A2 (.I(_03337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11130__B (.I(_03347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11131__I (.I(_03348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11133__A1 (.I(_03345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11133__A2 (.I(_03346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11133__B (.I(_03350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11135__A2 (.I(_03352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11138__A2 (.I(_03337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11145__B (.I(_03361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11146__I (.I(_03362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11148__A1 (.I(_03360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11148__B (.I(_03364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11150__A2 (.I(_03366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11153__A2 (.I(_03352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11161__I (.I(_03376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11162__I (.I(_03377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11165__B (.I(_03380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11166__I (.I(_03381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11168__A1 (.I(_03374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11168__A2 (.I(_03378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11168__B (.I(_03383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11170__A2 (.I(_03385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11173__A2 (.I(_03366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11180__I (.I(_03221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11182__B (.I(_03396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11184__A1 (.I(_03394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11184__A2 (.I(_03395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11184__B (.I(_03398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11187__A1 (.I(\filters.high[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11189__A2 (.I(_03403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11192__A2 (.I(_03385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11199__B (.I(_03412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11200__A1 (.I(_03411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11200__B (.I(_03413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11201__A1 (.I(_03410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11205__A2 (.I(_03403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11210__I (.I(\filters.band[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11211__I (.I(_03395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11213__A1 (.I(_03422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11216__A1 (.I(\filters.high[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11240__A1 (.I(_03243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11240__B1 (.I(_03245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11247__A2 (.I(_03226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11249__A1 (.I(_03236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11259__A1 (.I(_03468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11259__A2 (.I(_03226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11260__A1 (.I(_03202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11260__A2 (.I(_03194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11261__I (.I(_03470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11263__I (.I(_03472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11264__I (.I(_03473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11267__I (.I(_03476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11268__B (.I(_03236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11269__A2 (.I(_03236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11273__A1 (.I(_03243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11273__B1 (.I(_03245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11274__A1 (.I(_02088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11276__I (.I(_02334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11277__A1 (.I(\filters.cutoff_lut[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11278__A1 (.I(_02308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11279__A1 (.I(\filters.cutoff_lut[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11280__A1 (.I(_02314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11281__A1 (.I(\filters.cutoff_lut[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11282__A1 (.I(_02316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11284__I (.I(net14));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11287__A2 (.I(_01003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11288__A2 (.I(_01093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11289__A1 (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11289__A2 (.I(_03494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11293__I (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11295__A1 (.I(_03499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11296__C (.I(_02273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11298__A1 (.I(_02314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11299__I (.I(_02334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11301__A1 (.I(_02316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11303__A1 (.I(_02299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11305__A1 (.I(_01812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11306__I (.I(_03507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11307__I (.I(_03507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11308__A1 (.I(_03499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11309__C (.I(_02273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11310__I (.I(_02184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11312__A1 (.I(_03511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11313__I (.I(_02187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11315__A1 (.I(_03513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11319__B (.I(_03517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11320__A1 (.I(_03515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11326__A1 (.I(_01740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11328__A1 (.I(_02103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11329__B (.I(_03517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11330__A1 (.I(_03511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11331__B (.I(_03517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11332__A1 (.I(_03513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11333__B (.I(_03517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11334__A1 (.I(_03515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11335__S0 (.I(_01146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11335__S1 (.I(_01160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11336__I (.I(_03529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11337__S0 (.I(_01147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11337__S1 (.I(_01161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11338__A2 (.I(_03531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11339__I (.I(_03532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11342__I (.I(_02710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11343__A1 (.I(_02707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11343__A2 (.I(_02711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11344__A1 (.I(_03039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11349__A1 (.I(_03535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11350__A1 (.I(_02847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11351__A1 (.I(_01585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11351__A2 (.I(_03534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11351__A3 (.I(_03544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11352__A1 (.I(_03534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11352__A2 (.I(_03544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11353__A1 (.I(\channels.ctrl_reg2[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11353__A2 (.I(_01282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11354__A1 (.I(\channels.ctrl_reg3[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11354__A2 (.I(_01581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11354__B1 (.I(_01295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11354__B2 (.I(\channels.ctrl_reg1[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11356__A1 (.I(_03529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11356__A2 (.I(_03531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11357__A2 (.I(_03549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11358__A1 (.I(_01254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11361__A1 (.I(_01585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11361__A2 (.I(_03529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11361__A3 (.I(_03531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11361__A4 (.I(_03549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11367__B2 (.I(_03558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11368__I (.I(_02974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11370__A1 (.I(_03138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11372__B2 (.I(_03558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11374__A1 (.I(_03138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11376__B1 (.I(_01372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11376__B2 (.I(_03558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11378__A1 (.I(_03138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11380__B2 (.I(_03558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11383__A1 (.I(_03566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11385__I (.I(_01089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11386__I (.I(_01240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11387__B1 (.I(_01420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11388__I (.I(_02974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11390__A1 (.I(_03566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11392__B1 (.I(_01448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11394__A1 (.I(_03566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11396__B1 (.I(_01475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11398__A1 (.I(_03566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11400__B1 (.I(_01503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11403__A1 (.I(_03578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11405__I (.I(_01089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11406__I (.I(_01240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11407__B1 (.I(_01524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11408__A2 (.I(_01245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11408__B1 (.I(_01530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11411__B1 (.I(_01539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11413__A1 (.I(_03578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11415__B1 (.I(_01552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11417__A1 (.I(_03578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11418__B1 (.I(_01568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11420__A1 (.I(_03578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11425__B2 (.I(_03592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11426__I (.I(_03149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11427__A2 (.I(_03593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11430__B2 (.I(_03592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11431__A2 (.I(_03593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11434__B1 (.I(_01372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11434__B2 (.I(_03592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11435__A2 (.I(_03593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11438__B2 (.I(_03592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11439__I (.I(_02364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11440__A2 (.I(_03593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11441__A1 (.I(_03600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11443__I (.I(_01104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11444__I (.I(_01219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11445__B1 (.I(_01420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11446__I (.I(_03149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11447__A2 (.I(_03605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11448__A1 (.I(_03600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11450__B1 (.I(_01448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11451__A2 (.I(_03605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11452__A1 (.I(_03600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11454__B1 (.I(_01475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11455__A2 (.I(_03605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11456__A1 (.I(_03600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11458__B1 (.I(_01503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11459__I (.I(_02364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11460__A2 (.I(_03605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11461__A1 (.I(_03612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11463__I (.I(_01104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11464__I (.I(_01219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11465__B1 (.I(_01524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11466__A2 (.I(_01230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11466__B1 (.I(_01530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11469__B1 (.I(_01539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11471__A1 (.I(_03612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11473__B1 (.I(_01552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11475__A1 (.I(_03612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11476__B1 (.I(_01568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11478__A1 (.I(_03612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11481__I (.I(_00389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11482__A1 (.I(_02289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11482__A2 (.I(_01954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11483__I (.I(_03624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11484__I (.I(_03624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11486__A1 (.I(\channels.freq1[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11487__A1 (.I(_02308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11488__A1 (.I(\channels.freq1[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11489__A1 (.I(_03511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11490__A1 (.I(\channels.freq1[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11491__A1 (.I(_03513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11492__A1 (.I(\channels.freq1[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11493__A1 (.I(_03515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11494__I (.I(_03624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11495__I (.I(_03624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11497__A1 (.I(\channels.freq1[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11498__A1 (.I(_02319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11499__A1 (.I(\channels.freq1[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11500__A1 (.I(_02324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11501__A1 (.I(\channels.freq1[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11502__A1 (.I(_02326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11503__A1 (.I(\channels.freq1[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11504__A1 (.I(_02328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11505__I (.I(_01740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11506__I (.I(_01779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11508__I (.I(_03641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11509__I (.I(_03641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11511__A1 (.I(\channels.pw1[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11512__A1 (.I(_03639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11513__A1 (.I(\channels.pw1[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11514__A1 (.I(_03511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11515__A1 (.I(\channels.pw1[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11516__A1 (.I(_03513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11517__A1 (.I(\channels.pw1[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11518__A1 (.I(_03515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11519__I (.I(_03641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11520__I (.I(_03641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11523__A1 (.I(\channels.pw1[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11524__A1 (.I(_02319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11525__A1 (.I(\channels.pw1[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11526__A1 (.I(_02324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11527__A1 (.I(\channels.pw1[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11528__A1 (.I(_02326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11529__A1 (.I(\channels.pw1[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11530__A1 (.I(_02328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11536__A1 (.I(_03639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11537__I (.I(_01755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11539__A1 (.I(_03662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11541__A1 (.I(\channels.freq2[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11542__A1 (.I(_03664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11545__A1 (.I(_03666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11546__I (.I(_02149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11551__A1 (.I(_03668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11552__I (.I(_02154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11554__A1 (.I(_03673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11555__I (.I(_01812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11557__A1 (.I(_03675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11558__I (.I(_01817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11560__A1 (.I(_03677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11561__A2 (.I(_01871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11565__A1 (.I(\channels.freq3[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11566__A1 (.I(_03639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11567__A1 (.I(\channels.freq3[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11568__A1 (.I(_03662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11569__A1 (.I(\channels.freq3[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11570__A1 (.I(_03664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11571__A1 (.I(\channels.freq3[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11572__A1 (.I(_03666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11577__A1 (.I(\channels.freq3[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11578__A1 (.I(_03668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11580__A1 (.I(_03673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11582__A1 (.I(_03675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11583__A1 (.I(\channels.freq3[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11584__A1 (.I(_03677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11589__A1 (.I(\channels.pw3[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11590__A1 (.I(_03639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11591__A1 (.I(\channels.pw3[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11592__A1 (.I(_03662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11593__A1 (.I(\channels.pw3[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11594__A1 (.I(_03664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11595__A1 (.I(\channels.pw3[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11596__A1 (.I(_03666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11600__A1 (.I(\channels.pw3[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11601__A1 (.I(_03668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11602__A1 (.I(\channels.pw3[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11603__A1 (.I(_03673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11604__A1 (.I(\channels.pw3[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11605__A1 (.I(_03675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11607__A1 (.I(_03677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11608__I (.I(_01740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11609__A1 (.I(_01780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11610__I (.I(_03711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11611__I (.I(_03711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11613__A1 (.I(\channels.pw2[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11614__A1 (.I(_03710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11615__A1 (.I(\channels.pw2[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11616__A1 (.I(_03662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11617__A1 (.I(\channels.pw2[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11618__A1 (.I(_03664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11619__A1 (.I(\channels.pw2[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11620__A1 (.I(_03666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11621__I (.I(_03711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11622__I (.I(_03711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11624__I (.I(_03721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11625__A1 (.I(\channels.pw2[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11625__B (.I(_03722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11626__A1 (.I(_03668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11627__A1 (.I(\channels.pw2[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11627__B (.I(_03722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11628__A1 (.I(_03673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11629__B (.I(_03722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11630__A1 (.I(_03675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11631__B (.I(_03722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11632__A1 (.I(_03677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11633__A2 (.I(_01093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11636__I (.I(_03729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11637__I (.I(_03730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11638__I (.I(_03731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11639__I (.I(_01750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11640__I (.I(_03733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11642__A1 (.I(\channels.clk_div[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11642__B (.I(_03735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11643__A1 (.I(_03728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11645__A2 (.I(_03728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11647__A1 (.I(_02272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11650__A1 (.I(_01933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11651__I (.I(_02839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11653__I (.I(_01319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11654__I (.I(_03131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11655__I (.I(_03039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11656__I (.I(_02721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11657__I (.I(_02687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11663__A1 (.I(_03535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11665__A2 (.I(_03531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11667__A1 (.I(\channels.sus_rel1[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11668__A1 (.I(\channels.sus_rel3[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11668__B2 (.I(\channels.sus_rel2[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11669__A2 (.I(_03759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11670__A2 (.I(_03759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11671__A1 (.I(\channels.sus_rel1[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11672__A1 (.I(\channels.sus_rel3[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11672__B2 (.I(\channels.sus_rel2[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11673__I0 (.I(_02711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11673__S (.I(_03763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11674__A1 (.I(\channels.sus_rel3[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11675__A1 (.I(\channels.sus_rel2[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11675__B1 (.I(_01295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11675__B2 (.I(\channels.sus_rel1[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11676__A1 (.I(_01168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11677__A1 (.I(_01168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11678__A1 (.I(\channels.sus_rel3[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11679__A1 (.I(\channels.sus_rel2[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11679__B2 (.I(\channels.sus_rel1[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11681__B1 (.I(_03771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11682__A2 (.I(_02711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11682__B1 (.I(_03131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11682__B2 (.I(_03766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11683__A2 (.I(_02752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11683__B1 (.I(_03766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11683__B2 (.I(_03039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11684__A2 (.I(_03535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11685__A1 (.I(_03535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11685__A2 (.I(_03771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11687__A2 (.I(_03755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11687__B1 (.I(_03757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11687__B2 (.I(_03777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11688__A1 (.I(_03534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11690__A1 (.I(\channels.sus_rel3[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11690__B2 (.I(\channels.sus_rel2[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11694__I (.I(_03784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11695__B2 (.I(\channels.atk_dec2[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11696__A1 (.I(_03757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11698__I0 (.I(\channels.atk_dec1[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11698__S (.I(_03784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11699__A2 (.I(_03789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11700__I (.I(_03532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11701__B2 (.I(\channels.atk_dec2[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11701__C2 (.I(\channels.atk_dec1[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11704__B2 (.I(\channels.atk_dec2[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11705__A1 (.I(\channels.sus_rel3[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11705__B2 (.I(\channels.sus_rel2[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11707__I0 (.I(\channels.atk_dec1[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11707__S (.I(_03784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11708__A2 (.I(_03798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11708__B (.I(_03532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11709__B2 (.I(\channels.atk_dec2[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11709__C2 (.I(\channels.atk_dec1[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11715__A1 (.I(\channels.sus_rel3[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11715__B2 (.I(\channels.sus_rel2[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11716__A1 (.I(\channels.atk_dec3[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11716__B2 (.I(\channels.atk_dec2[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11717__A1 (.I(_03757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11718__I0 (.I(\channels.atk_dec1[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11718__I1 (.I(\channels.sus_rel1[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11718__S (.I(_03784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11719__A2 (.I(_03809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11720__B2 (.I(\channels.atk_dec2[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11720__C2 (.I(\channels.atk_dec1[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11726__A1 (.I(\channels.atk_dec3[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11726__B2 (.I(\channels.atk_dec2[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11727__A1 (.I(\channels.sus_rel3[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11727__B2 (.I(\channels.sus_rel2[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11728__S (.I(_03757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11729__I0 (.I(\channels.atk_dec1[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11729__I1 (.I(\channels.sus_rel1[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11731__B2 (.I(\channels.atk_dec2[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11731__C2 (.I(\channels.atk_dec1[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11740__I (.I(_01150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11742__S0 (.I(_03832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11742__S1 (.I(_01171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11751__I (.I(_01166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11752__S0 (.I(_03832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11752__S1 (.I(_03842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11763__S0 (.I(_03832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11763__S1 (.I(_03842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11770__S0 (.I(_01152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11770__S1 (.I(_01171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11775__S1 (.I(_01167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11783__S1 (.I(_01167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11784__A2 (.I(_03874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11788__S0 (.I(_01151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11788__S1 (.I(_01167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11792__A2 (.I(_03874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11795__I (.I(_01149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11796__S0 (.I(_03886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11796__S1 (.I(_01166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11797__I (.I(_03887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11801__S0 (.I(_03886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11801__S1 (.I(_01170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11802__A3 (.I(_03887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11807__S0 (.I(_01150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11807__S1 (.I(_01165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11812__S0 (.I(_01151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11812__S1 (.I(_03842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11813__A2 (.I(_03903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11814__S0 (.I(_03832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11814__S1 (.I(_01171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11817__A1 (.I(_03905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11818__S0 (.I(_01150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11818__S1 (.I(_01166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11823__I (.I(_03905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11825__S (.I(_03886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11828__A1 (.I(_01151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11828__C (.I(_01170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11829__A1 (.I(_03842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11834__S0 (.I(_03886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11834__S1 (.I(_01170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11835__A2 (.I(_03925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11836__A2 (.I(_03925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11838__A1 (.I(_01584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11839__A2 (.I(_03903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11844__I (.I(_03934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11845__A2 (.I(_03935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11846__I (.I(_03936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11847__A1 (.I(_03744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11850__A1 (.I(_03744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11850__B (.I(_03940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11855__A2 (.I(_03934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11856__I (.I(_03945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11862__I (.I(_03945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11880__A2 (.I(_03964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11882__A1 (.I(_02752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11890__A2 (.I(_03974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11893__A1 (.I(_03128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11895__A2 (.I(_03978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11903__A1 (.I(_03905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11912__A1 (.I(_01584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11920__A1 (.I(_03534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11920__A2 (.I(_04002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11920__B (.I(_01585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11921__A1 (.I(_04001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11923__A1 (.I(_02356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11924__I (.I(_04006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11926__I (.I(_03935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11928__A1 (.I(_01581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11928__B (.I(_01102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11929__I (.I(_04011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11933__A2 (.I(_03874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11934__A2 (.I(_03874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11938__I (.I(_04001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11940__A1 (.I(_04019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11948__I (.I(_04006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11950__A1 (.I(_04019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11951__I (.I(_04011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11960__A1 (.I(_04019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11963__A1 (.I(_03903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11964__B (.I(_03903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11965__A1 (.I(_03935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11968__I (.I(_04006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11969__I (.I(_04001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11972__A1 (.I(_04044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11973__I (.I(_04011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11977__A1 (.I(_04019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11983__A1 (.I(_04044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11989__A1 (.I(_04001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11993__A1 (.I(_04044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11998__A1 (.I(_04044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12002__A1 (.I(_03925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12002__B (.I(_03935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12003__A1 (.I(_03925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12006__A1 (.I(_02363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12007__I (.I(_04074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12009__B (.I(_01032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12010__I (.I(_04077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12020__I (.I(_04074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12021__I (.I(_04077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12030__I (.I(_04074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12031__I (.I(_04077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12050__A2 (.I(_02354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12053__A1 (.I(_04101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12054__A1 (.I(_03744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12055__I (.I(_04103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12057__A1 (.I(_01319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12057__B (.I(_01032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12058__I (.I(_04106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12068__I (.I(_04103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12069__I (.I(_04106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12078__I (.I(_04103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12079__I (.I(_04106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12094__A1 (.I(_01240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12099__A1 (.I(_01219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12152__I (.I(_01093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12153__A1 (.I(_04158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12153__A2 (.I(_03226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12154__I (.I(_04159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12155__I (.I(_04160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12156__A4 (.I(\filters.high[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12158__I (.I(_04163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12159__A1 (.I(_03317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12165__A1 (.I(\filters.res_lut[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12165__A2 (.I(_04170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12166__A2 (.I(_04171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12167__A1 (.I(\filters.res_lut[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12168__I (.I(_04173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12171__A4 (.I(\filters.high[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12172__A2 (.I(_04177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12177__A1 (.I(_04176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12177__A2 (.I(_04182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12178__A1 (.I(\filters.res_lut[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12179__I (.I(_04184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12180__I (.I(_04185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12181__I (.I(_04186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12184__A1 (.I(_03239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12184__A3 (.I(_04189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12185__I (.I(_04190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12187__A1 (.I(_03350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12187__A3 (.I(_04192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12188__A4 (.I(\filters.high[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12192__A1 (.I(\filters.res_lut[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12193__I (.I(_04198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12194__I (.I(_04199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12195__I (.I(_04200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12196__A1 (.I(_03288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12200__I (.I(_04182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12201__A1 (.I(\filters.res_lut[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12202__I (.I(_04207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12206__A3 (.I(_04211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12207__A2 (.I(_04210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12207__B (.I(_04212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12209__A1 (.I(_03239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12209__A3 (.I(_04189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12210__I (.I(_04215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12212__I0 (.I(\filters.cutoff_lut[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12213__I (.I(_04218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12214__I (.I(_04219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12215__I (.I(_04220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12216__I (.I(_04221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12217__A1 (.I(_03200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12217__A3 (.I(_04222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12218__A4 (.I(\filters.high[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12221__A1 (.I(\filters.res_lut[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12222__I (.I(_04227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12224__I (.I(_04229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12226__A3 (.I(_04231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12228__A3 (.I(_04221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12229__I0 (.I(\filters.cutoff_lut[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12230__I (.I(_04235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12233__A1 (.I(_03200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12233__A3 (.I(_04238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12234__A4 (.I(\filters.high[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12238__A1 (.I(_03273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12238__A3 (.I(_04231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12240__A1 (.I(_04233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12240__A2 (.I(_04245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12242__A1 (.I(_04233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12242__A2 (.I(_04245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12247__I (.I(_04235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12249__I (.I(_04254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12250__A3 (.I(_04255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12251__I (.I(_04218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12252__I (.I(_04257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12253__I (.I(_04258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12254__A3 (.I(_04259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12255__A1 (.I(_03288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12256__A1 (.I(\filters.res_lut[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12257__A1 (.I(_04261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12260__I (.I(_04265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12261__A1 (.I(_03348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12261__A2 (.I(_04190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12264__A1 (.I(_04266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12264__A2 (.I(_04269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12266__A1 (.I(_03362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12266__A2 (.I(_04271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12269__A1 (.I(_04274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12273__I (.I(_04278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12276__A1 (.I(_04281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12278__A1 (.I(_04252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12278__A3 (.I(_04283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12280__A1 (.I(\filters.res_lut[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12281__I (.I(_04286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12286__I (.I(_04291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12288__I (.I(_04198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12290__I (.I(_04295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12291__I (.I(_04281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12292__B1 (.I(_04296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12292__B2 (.I(_04297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12293__A1 (.I(_04281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12293__A2 (.I(_04291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12293__A4 (.I(_04296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12295__I (.I(_04269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12296__I (.I(_04207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12305__A1 (.I(_03199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12306__I (.I(_04311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12308__I0 (.I(\filters.cutoff_lut[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12309__I (.I(_04314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12310__I (.I(_04315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12311__I (.I(_04316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12313__A2 (.I(_04318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12317__I0 (.I(\filters.cutoff_lut[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12317__I1 (.I(\filters.res_lut[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12318__I (.I(_04323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12319__I (.I(_04324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12321__A1 (.I(_04322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12321__A2 (.I(_04326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12322__A1 (.I(_04319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12322__A2 (.I(_04327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12327__A1 (.I(_03302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12327__A2 (.I(_04332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12330__A2 (.I(_04219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12334__A1 (.I(_04291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12334__A2 (.I(_04266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12336__I (.I(_04341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12337__A1 (.I(_03383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12337__A3 (.I(_04185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12338__A1 (.I(_03316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12338__A3 (.I(_04199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12343__A1 (.I(_04252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12344__A1 (.I(_04252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12345__A2 (.I(_04283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12350__A2 (.I(_04355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12351__A1 (.I(_04252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12351__A3 (.I(_04283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12353__A1 (.I(_04356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12359__A1 (.I(_04319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12359__A2 (.I(_04327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12360__I (.I(_04323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12361__I (.I(_04366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12362__A2 (.I(_03270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12364__A1 (.I(_04367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12364__A2 (.I(_04369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12365__I (.I(_04314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12366__I (.I(_04371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12367__A1 (.I(_04372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12368__I0 (.I(\filters.cutoff_lut[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12370__I (.I(_04375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12371__I (.I(_04376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12372__I (.I(_04377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12373__A2 (.I(_04378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12375__A2 (.I(_04380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12381__A1 (.I(_04229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12385__A2 (.I(_04390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12386__I (.I(_04258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12387__A1 (.I(_04392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12389__A1 (.I(_03381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12389__A2 (.I(_04341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12390__I (.I(_04395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12392__A1 (.I(_04265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12392__A2 (.I(_04397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12393__A1 (.I(_04200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12394__I (.I(_04184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12395__I (.I(_04400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12396__A4 (.I(\filters.high[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12398__A1 (.I(_03398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12398__A2 (.I(_04403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12401__A1 (.I(_04401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12401__A2 (.I(_04406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12411__A2 (.I(_04416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12415__A2 (.I(_04420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12437__A1 (.I(\filters.cutoff_lut[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12439__I (.I(_04444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12441__I (.I(_04446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12442__A2 (.I(_04447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12443__I (.I(_04372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12444__I (.I(_04375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12445__I (.I(_04450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12446__I (.I(_04451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12447__I (.I(_04452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12448__A2 (.I(_04322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12448__B1 (.I(_04453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12449__A4 (.I(_04453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12451__A1 (.I(_04366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12451__A2 (.I(_04390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12452__A3 (.I(_04376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12453__A1 (.I(_03273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12453__A2 (.I(_04372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12454__A2 (.I(_04458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12454__A3 (.I(_04459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12455__A1 (.I(_04456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12456__A1 (.I(_04448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12460__A1 (.I(_04319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12460__A2 (.I(_04327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12460__A3 (.I(_04380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12461__I (.I(_04254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12462__I (.I(_04390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12464__I (.I(_04257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12466__A2 (.I(_04468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12466__B2 (.I(_04471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12468__A2 (.I(_04471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12468__A3 (.I(_04390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12470__I (.I(_04227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12472__A2 (.I(_04476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12473__A2 (.I(_04278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12475__A1 (.I(_04220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12475__A2 (.I(_04480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12480__A1 (.I(_04199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12481__I (.I(_04185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12482__A4 (.I(_03410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12483__A1 (.I(_03413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12483__A2 (.I(_04488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12484__I (.I(_04489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12486__A1 (.I(_04487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12488__A1 (.I(_04475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12488__A2 (.I(_04482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12492__I (.I(_04416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12493__A2 (.I(_04498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12495__A2 (.I(_04500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12499__I (.I(_04406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12501__A1 (.I(_04504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12501__B2 (.I(_04506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12502__A2 (.I(_04504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12502__A3 (.I(_04182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12507__A1 (.I(_04512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12517__A1 (.I(_03333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12518__A1 (.I(_03273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12518__A3 (.I(_04296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12519__I (.I(_04266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12520__A1 (.I(_03317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12520__A2 (.I(_04525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12524__A1 (.I(_03333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12524__A2 (.I(_04529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12526__A1 (.I(_04233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12526__A2 (.I(_04245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12527__A2 (.I(_04528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12528__A2 (.I(_04210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12530__A1 (.I(_04535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12530__A2 (.I(_04171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12531__A1 (.I(\filters.res_lut[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12534__A1 (.I(_04537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12535__A1 (.I(\filters.res_lut[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12536__A2 (.I(_04541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12540__A2 (.I(_04210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12543__A1 (.I(_04356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12554__A1 (.I(_04528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12555__I (.I(_04500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12556__I (.I(_04561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12557__A1 (.I(_04468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12557__A2 (.I(_04562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12558__A1 (.I(_04535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12558__A2 (.I(_04537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12559__A1 (.I(_03317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12559__A2 (.I(_04506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12561__A2 (.I(_04566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12561__A3 (.I(_04504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12565__A1 (.I(_04297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12565__A2 (.I(_04498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12569__I (.I(_04231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12571__A2 (.I(_04576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12572__I (.I(_04525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12573__A1 (.I(_03302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12573__A2 (.I(_04332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12573__A3 (.I(_04578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12579__A1 (.I(_04583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12580__A1 (.I(_04574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12582__A1 (.I(_04574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12583__A1 (.I(_04583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12588__I (.I(_04593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12589__A2 (.I(_04171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12590__I (.I(_04529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12591__I (.I(_04596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12592__A1 (.I(_04468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12592__A2 (.I(_04597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12593__I (.I(_04506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12594__I (.I(_04296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12596__A1 (.I(_04297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12596__B1 (.I(_04601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12597__A2 (.I(_04297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12597__A4 (.I(_04601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12599__A1 (.I(_04261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12599__A2 (.I(_04541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12607__A1 (.I(_03256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12607__A2 (.I(_04566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12608__A2 (.I(_04171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12609__I (.I(_04369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12610__I (.I(_04578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12612__A2 (.I(_04468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12612__A3 (.I(_04616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12612__A4 (.I(_04617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12613__I (.I(_04498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12614__A2 (.I(_04619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12616__A1 (.I(_04541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12623__I (.I(_04420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12625__I (.I(_04630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12626__I (.I(_04619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12627__I (.I(_04616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12628__I (.I(_04617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12629__A1 (.I(_03256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12629__A2 (.I(_04566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12630__A2 (.I(_04632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12631__A1 (.I(_03256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12631__A2 (.I(_04566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12632__A2 (.I(_04541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12633__A2 (.I(_04631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12634__A2 (.I(_04631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12635__I (.I(_04207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12636__I (.I(_04641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12637__I (.I(_04642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12639__I (.I(_04644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12640__A2 (.I(_04645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12642__A1 (.I(\filters.res_lut[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12642__A2 (.I(_04170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12643__A2 (.I(_04537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12643__B2 (.I(_04261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12647__A1 (.I(_04535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12648__A2 (.I(_04601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12650__I0 (.I(_04644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12659__A1 (.I(_04322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12661__I (.I(_04632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12662__A1 (.I(_04667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12672__A1 (.I(_04674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12672__A2 (.I(_04675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12676__A2 (.I(_04674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12676__A3 (.I(_04675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12676__B (.I(_04681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12691__I (.I(_04392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12692__A1 (.I(_04694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12692__A2 (.I(_04281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12692__B2 (.I(_04697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12693__I (.I(_04255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12694__A1 (.I(_04699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12694__A2 (.I(_04697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12696__A2 (.I(_04480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12697__I (.I(_04257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12699__I (.I(_04476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12700__A1 (.I(_04705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12702__A1 (.I(_04701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12703__A1 (.I(_04265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12704__I (.I(_03184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12705__I0 (.I(\filters.high[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12705__I1 (.I(\filters.band[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12705__S (.I(_04710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12706__I (.I(_04711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12707__I (.I(_04712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12708__A1 (.I(_04186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12708__A2 (.I(_04713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12709__A1 (.I(_04274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12709__A2 (.I(_04295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12710__A2 (.I(_04714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12712__A1 (.I(_04701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12714__A1 (.I(_04366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12715__A3 (.I(_04376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12716__A1 (.I(_03288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12716__A2 (.I(_04316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12718__A1 (.I(_04458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12718__A2 (.I(_04459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12719__A1 (.I(_04458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12719__A2 (.I(_04459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12724__A1 (.I(_04728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12724__B2 (.I(_04259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12725__A1 (.I(_04728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12725__A2 (.I(_04259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12729__A1 (.I(_04258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12731__I (.I(_04711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12732__A1 (.I(_04173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12732__A2 (.I(_04737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12733__S (.I(_04710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12734__I (.I(_04739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12735__A1 (.I(_04184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12735__A2 (.I(_04740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12736__I (.I(_04198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12737__A2 (.I(_04742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12738__A3 (.I(_04743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12739__A1 (.I(_04732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12744__I (.I(_04489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12745__I (.I(_04750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12746__I (.I(_04751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12748__A1 (.I(_04286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12748__A2 (.I(_04753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12749__A2 (.I(_04743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12750__A2 (.I(_04743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12752__I (.I(_04713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12753__I (.I(_04758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12754__A1 (.I(_04641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12758__I (.I(_04211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12759__I (.I(_04764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12760__I (.I(_04753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12761__A1 (.I(_04714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12762__A1 (.I(_04714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12764__A2 (.I(_04766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12765__A2 (.I(_04766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12771__A1 (.I(\filters.cutoff_lut[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12771__A2 (.I(_04776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12772__A1 (.I(_04593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12773__A1 (.I(\filters.cutoff_lut[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12775__I (.I(_04780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12776__A1 (.I(_03200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12776__A3 (.I(_04781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12777__A1 (.I(\filters.cutoff_lut[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12778__I (.I(_04783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12779__A3 (.I(_04784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12785__I (.I(_04783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12786__A1 (.I(_04311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12786__A3 (.I(_04444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12787__A2 (.I(_04323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12789__A2 (.I(_04314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12791__A1 (.I(_04792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12791__A2 (.I(_04796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12793__A1 (.I(_04787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12795__I (.I(_04800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12797__I (.I(_04783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12798__I (.I(_04803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12799__I (.I(_04804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12800__I (.I(_04805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12801__A1 (.I(_04322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12801__A2 (.I(_04802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12801__B1 (.I(_04806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12802__A1 (.I(_04792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12802__A2 (.I(_04807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12809__A1 (.I(_04787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12810__A1 (.I(\filters.cutoff_lut[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12813__I (.I(_04818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12816__A3 (.I(_04444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12817__A3 (.I(_04784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12818__I (.I(_04780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12820__A3 (.I(_04825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12822__A1 (.I(_04821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12822__A2 (.I(_04827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12828__A1 (.I(_04324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12829__A1 (.I(_04316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12829__A2 (.I(_04480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12830__A2 (.I(_04377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12832__A1 (.I(_04831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12832__A2 (.I(_04833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12832__A3 (.I(_04837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12835__A1 (.I(_04732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12837__A1 (.I(_04732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12839__A1 (.I(_04792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12839__A2 (.I(_04796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12841__I (.I(_04220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12843__A1 (.I(_04847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12843__A2 (.I(_04269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12843__B2 (.I(_04848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12845__A1 (.I(_04848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12845__A2 (.I(_04850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12847__A1 (.I(_04476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12848__I (.I(_04271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12849__A1 (.I(_03364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12849__A2 (.I(_04219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12850__A3 (.I(_04192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12851__A1 (.I(_04853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12851__A2 (.I(_04855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12851__A3 (.I(_04856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12852__I (.I(_04739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12853__A2 (.I(_04858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12854__S (.I(_04710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12855__I (.I(_04860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12857__A1 (.I(_04400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12859__A1 (.I(_04200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12859__A2 (.I(_04864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12860__A2 (.I(_04863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12861__A1 (.I(_04852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12862__A2 (.I(_04846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12863__A2 (.I(_04844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12872__A1 (.I(_04821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12872__A2 (.I(_04827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12873__A1 (.I(\filters.cutoff_lut[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12877__A1 (.I(_03199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12877__A2 (.I(_04215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12879__A3 (.I(_04884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12881__A1 (.I(_03302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12881__A2 (.I(_04332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12881__A3 (.I(_04800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12882__A3 (.I(_04803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12885__A1 (.I(_04886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12885__A2 (.I(_04890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12886__B1 (.I(_04378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12887__I (.I(_04316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12888__A1 (.I(_04893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12888__A4 (.I(_04378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12891__A1 (.I(_04261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12891__A2 (.I(_04896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12895__A1 (.I(_04367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12896__A2 (.I(_04371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12897__A1 (.I(_03316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12897__A2 (.I(_04163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12897__A3 (.I(_04450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12898__A1 (.I(_04902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12898__A2 (.I(_04903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12900__A1 (.I(_04895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12900__A2 (.I(_04900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12900__A3 (.I(_04905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12902__A1 (.I(_04852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12904__A1 (.I(_04852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12906__A1 (.I(_04833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12906__A2 (.I(_04837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12907__A1 (.I(_04833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12907__A2 (.I(_04837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12908__A1 (.I(_04831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12909__A1 (.I(_04855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12909__A2 (.I(_04856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12910__A1 (.I(_04855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12910__A2 (.I(_04856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12911__A1 (.I(_04853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12912__A1 (.I(_04229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12916__A1 (.I(_04921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12919__A2 (.I(_04924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12920__S (.I(_03185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12921__I (.I(_04926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12922__A1 (.I(_04487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12922__A2 (.I(_04927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12924__A1 (.I(_04295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12924__A2 (.I(_04929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12925__A2 (.I(_04928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12930__A1 (.I(_04632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12931__A1 (.I(_04644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12933__A1 (.I(_04846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12934__A1 (.I(_04844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12936__A1 (.I(_04863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12937__A1 (.I(_04863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12939__I (.I(_04858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12941__A1 (.I(_04416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12941__A2 (.I(_04946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12944__A1 (.I(_04938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12947__A1 (.I(_04475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12947__A2 (.I(_04482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12949__A1 (.I(_04475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12949__A2 (.I(_04482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12951__A1 (.I(_04456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12952__A1 (.I(_04701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12956__A2 (.I(_04766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12959__A1 (.I(_04512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12959__A2 (.I(_04420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12964__A1 (.I(_04619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12964__A2 (.I(_04966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12965__A1 (.I(_04619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12965__A2 (.I(_04966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12970__A1 (.I(_04448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12986__A1 (.I(_04952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12986__A2 (.I(_04991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12988__A1 (.I(_04512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12988__A2 (.I(_04642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12993__A1 (.I(_04211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12993__A2 (.I(_04966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12995__A2 (.I(_05000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12997__A2 (.I(_05000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12998__A1 (.I(_04996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13003__A1 (.I(_04996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13010__A1 (.I(_04993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13020__A1 (.I(_04996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13020__A3 (.I(_05000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13030__A1 (.I(_05035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13031__A2 (.I(_04992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13037__A1 (.I(_04992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13038__A1 (.I(_04952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13038__A2 (.I(_04991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13041__A1 (.I(_04952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13041__A2 (.I(_04991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13041__C (.I(_04993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13044__A1 (.I(_04928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13045__A1 (.I(_04928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13047__A2 (.I(_05049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13048__I (.I(_04946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13049__A1 (.I(_04641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13049__A2 (.I(_05049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13053__A2 (.I(_04921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13055__A1 (.I(_04900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13055__A2 (.I(_04905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13056__A1 (.I(_04900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13056__A2 (.I(_04905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13057__A1 (.I(_04895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13058__A1 (.I(_04699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13058__A2 (.I(_04291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13058__B2 (.I(_04697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13059__A1 (.I(_04699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13059__A2 (.I(_04221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13059__A3 (.I(_04274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13061__A1 (.I(_04705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13061__A2 (.I(_04751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13062__A1 (.I(_03398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13062__A2 (.I(_04219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13062__A3 (.I(_04403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13064__A2 (.I(_05069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13064__A3 (.I(_04341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13065__A2 (.I(_05070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13067__A1 (.I(_05066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13068__I (.I(_04926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13069__I (.I(_05074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13070__A2 (.I(_05075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13071__I1 (.I(\filters.band[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13071__S (.I(_03185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13072__I (.I(_05077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13073__I (.I(_05078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13074__A1 (.I(_04401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13075__A2 (.I(_04758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13076__A2 (.I(_05080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13081__A2 (.I(_05049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13082__A1 (.I(_05080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13083__A1 (.I(_05080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13085__I (.I(_04927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13087__A1 (.I(_04764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13087__A2 (.I(_05092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13096__A1 (.I(_04886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13096__A2 (.I(_04890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13098__A1 (.I(_03270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13100__A1 (.I(\filters.cutoff_lut[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13101__I (.I(_05106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13102__A1 (.I(_03199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13102__A2 (.I(_04215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13104__A2 (.I(_04163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13106__A2 (.I(_04332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13106__A3 (.I(_04783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13109__A2 (.I(_05114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13110__A1 (.I(_04902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13110__A2 (.I(_04903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13112__A1 (.I(_04535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13112__A2 (.I(_04896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13116__A1 (.I(_04367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13117__A2 (.I(_04315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13118__A3 (.I(_04450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13119__A2 (.I(_05124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13120__A1 (.I(_05122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13121__A2 (.I(_05121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13127__A2 (.I(_05114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13133__A1 (.I(_04369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13133__A2 (.I(_04818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13140__A2 (.I(_05145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13142__A2 (.I(_04800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13143__A1 (.I(_04278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13143__A2 (.I(_04780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13146__A1 (.I(_05142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13146__A2 (.I(_05147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13147__A2 (.I(_05124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13148__A1 (.I(_05122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13151__A2 (.I(_04896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13152__I (.I(_04366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13153__A1 (.I(_05158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13154__A1 (.I(_03348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13154__A3 (.I(_04375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13155__A2 (.I(_04315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13155__A3 (.I(_04271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13158__A2 (.I(_05157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13159__A1 (.I(_05138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13161__A1 (.I(_05066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13163__A1 (.I(_05121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13164__A1 (.I(_05121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13166__A2 (.I(_05070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13168__A2 (.I(_04737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13169__A1 (.I(_05069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13174__A1 (.I(\filters.band[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13174__A2 (.I(_05179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13175__A2 (.I(_03470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13176__A1 (.I(_05181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13176__A2 (.I(_04537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13177__I (.I(_04858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13178__A1 (.I(_04742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13180__I (.I(_05185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13182__A1 (.I(_04401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13182__A2 (.I(_05187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13183__A1 (.I(_05182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13183__A2 (.I(_05184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13183__A3 (.I(_05188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13193__A1 (.I(_05138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13195__A2 (.I(_05157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13196__A1 (.I(_05138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13198__A1 (.I(_05142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13198__A2 (.I(_05147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13199__I (.I(_05151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13200__A1 (.I(_05142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13200__A2 (.I(_05147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13203__A1 (.I(_04369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13203__B1 (.I(_05208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13204__A4 (.I(_05145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13208__A1 (.I(_03270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13208__A3 (.I(_05106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13211__A1 (.I(_05211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13211__A2 (.I(_05216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13212__A2 (.I(_04444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13214__I (.I(_04780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13215__A2 (.I(_05220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13224__I (.I(_04784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13226__A2 (.I(_05229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13227__A3 (.I(_04825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13229__A1 (.I(_04324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13230__A2 (.I(_04271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13230__A3 (.I(_04450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13231__A2 (.I(_04371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13232__A2 (.I(_05237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13234__A2 (.I(_05234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13239__A1 (.I(_05157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13240__A1 (.I(_05157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13242__A1 (.I(_04255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13242__A2 (.I(_04864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13242__B2 (.I(_04471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13243__A1 (.I(_04255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13243__A2 (.I(_04392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13243__A4 (.I(_04751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13245__A2 (.I(_04740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13246__A1 (.I(_05069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13246__A2 (.I(_04750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13247__A2 (.I(_04712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13249__A2 (.I(_05254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13251__A1 (.I(_04266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13252__A1 (.I(_04199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13253__I1 (.I(\filters.band[18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13253__S (.I(_03185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13254__I (.I(_05259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13255__A1 (.I(_04185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13255__A2 (.I(_05260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13258__A2 (.I(_05263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13262__I (.I(_05092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13263__A2 (.I(_05268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13264__A2 (.I(_05268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13269__A2 (.I(_05268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13270__A1 (.I(_05184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13270__A2 (.I(_05188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13271__A1 (.I(_05184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13271__A2 (.I(_05188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13273__I (.I(_05077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13276__A2 (.I(_05281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13298__A1 (.I(_05211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13298__A2 (.I(_05216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13304__A3 (.I(_05106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13308__A2 (.I(_04800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13309__A3 (.I(_04781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13309__A4 (.I(_04803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13310__A2 (.I(_04781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13310__B1 (.I(_04784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13314__A1 (.I(_05313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13317__A2 (.I(_05237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13318__A3 (.I(_05220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13318__A4 (.I(_04804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13319__B (.I(_05324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13320__A1 (.I(_04323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13320__A2 (.I(_04489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13321__A1 (.I(_04395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13321__A2 (.I(_04375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13322__A1 (.I(_04315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13328__A2 (.I(_05263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13329__A2 (.I(_05254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13330__A1 (.I(_05234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13331__A1 (.I(_05234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13333__B1 (.I(_04712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13334__A1 (.I(_04254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13334__A4 (.I(_04712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13336__A1 (.I(_04227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13336__A2 (.I(_04860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13337__A2 (.I(_04711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13338__A1 (.I(_04257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13338__A2 (.I(_04739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13340__A1 (.I(_05341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13340__A2 (.I(_05345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13341__I (.I(_05259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13342__A1 (.I(_04265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13343__A1 (.I(_04198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13343__A2 (.I(_04926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13344__S (.I(_04710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13345__I (.I(_05350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13346__A1 (.I(_04184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13349__A2 (.I(_05354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13353__A1 (.I(_04500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13353__A2 (.I(_05092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13359__A1 (.I(_04420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13359__A2 (.I(_05281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13361__I (.I(_05187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13362__A1 (.I(_04596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13365__A1 (.I(_04641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13367__A2 (.I(_05372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13372__A1 (.I(_05289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13372__A2 (.I(_05377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13398__A1 (.I(_05403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13398__A2 (.I(_05379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13402__A1 (.I(_04938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13410__A1 (.I(_05405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13410__A2 (.I(_05415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13415__A1 (.I(_05417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13415__A2 (.I(_05420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13418__A1 (.I(_05289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13418__A2 (.I(_05377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13419__A1 (.I(_05379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13419__A2 (.I(_05403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13421__A1 (.I(_05405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13421__A2 (.I(_05415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13422__A1 (.I(_05405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13422__A2 (.I(_05415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13422__B1 (.I(_05417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13422__B2 (.I(_05420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13424__A1 (.I(_05289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13424__A2 (.I(_05377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13426__A1 (.I(_05423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13426__A2 (.I(_05431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13434__I (.I(_04562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13435__A1 (.I(_05440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13435__A2 (.I(_05281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13435__A3 (.I(_05372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13439__A1 (.I(_04561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13440__I (.I(_04596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13441__I (.I(_05260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13444__A1 (.I(_05446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13446__A1 (.I(_04642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13447__A1 (.I(_05451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13449__A1 (.I(_05444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13449__A2 (.I(_05454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13459__I (.I(_05229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13460__I (.I(_04805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13461__A1 (.I(_04269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13461__A2 (.I(_04182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13463__I (.I(_04737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13464__A1 (.I(_05158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13464__A2 (.I(_05469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13465__A1 (.I(_04451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13471__A1 (.I(_05313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13471__B (.I(_05476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13473__A1 (.I(_03350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13473__A2 (.I(_04192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13473__A3 (.I(_05220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13474__A1 (.I(_03364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13474__A3 (.I(_04804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13479__A2 (.I(_04884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13480__A1 (.I(_04278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13480__A2 (.I(_05208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13482__A1 (.I(_04480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13482__A2 (.I(_05487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13484__A1 (.I(_05484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13484__A2 (.I(_05489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13489__I (.I(_05341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13490__A2 (.I(_05345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13491__A2 (.I(_05354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13492__A1 (.I(_05324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13496__A1 (.I(_04525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13497__A1 (.I(_04295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13499__I (.I(_05504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13500__A1 (.I(_04401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13503__I (.I(_04848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13504__I (.I(_04850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13505__A1 (.I(_05509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13505__A2 (.I(_04758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13505__B1 (.I(_04946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13505__B2 (.I(_05510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13507__A1 (.I(_05512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13507__A2 (.I(_05510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13507__A3 (.I(_04758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13507__A4 (.I(_04946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13509__A1 (.I(_04705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13509__A2 (.I(_05074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13510__I (.I(_04740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13511__A2 (.I(_05516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13513__A1 (.I(_04850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13515__A1 (.I(_05514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13515__A2 (.I(_05520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13516__A1 (.I(_05508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13525__A1 (.I(_05527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13525__A2 (.I(_05530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13529__A1 (.I(_05534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13529__A2 (.I(_03346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13534__I (.I(_04159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13535__I (.I(_03721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13538__A1 (.I(_03730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13539__I (.I(_05543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13540__I (.I(_05544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13541__I (.I(_05543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13542__I (.I(_05546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13544__A1 (.I(_05527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13544__A2 (.I(_05530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13549__A1 (.I(_05444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13549__A2 (.I(_05454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13555__I (.I(_04645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13557__A1 (.I(_05560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13557__A3 (.I(_05451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13558__I (.I(_04562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13559__A1 (.I(_05563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13564__A1 (.I(_04630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13566__A1 (.I(_04597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13566__A2 (.I(_05570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13568__A1 (.I(_04764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13568__A2 (.I(_05570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13571__A1 (.I(_05568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13575__I (.I(_05514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13576__A2 (.I(_05520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13577__A1 (.I(_05508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13580__I (.I(_05504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13581__A1 (.I(_04176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13583__I1 (.I(\filters.band[21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13583__S (.I(_05179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13584__A1 (.I(_04400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13584__A2 (.I(_05588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13587__A1 (.I(_04238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13587__B2 (.I(_04847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13588__A1 (.I(_04848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13588__A2 (.I(_04850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13590__A1 (.I(_04476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13590__A2 (.I(_05077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13592__A1 (.I(_04220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13592__A2 (.I(_04926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13593__A2 (.I(_05596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13593__A3 (.I(_05597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13594__A1 (.I(_05594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13595__A1 (.I(_05591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13596__A1 (.I(_05584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13606__A1 (.I(_05158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13606__A2 (.I(_05516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13607__A1 (.I(_04377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13607__A2 (.I(_04751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13608__A2 (.I(_04713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13612__A1 (.I(_05484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13612__A2 (.I(_05489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13614__A1 (.I(_04864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13615__A1 (.I(_03364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13615__A3 (.I(_05220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13616__A1 (.I(_03383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13616__A3 (.I(_04804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13617__A2 (.I(_05621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13619__I (.I(_05487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13620__I (.I(_05145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13622__A2 (.I(_05624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13622__B1 (.I(_05626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13623__A3 (.I(_05624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13623__A4 (.I(_05626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13625__A2 (.I(_04884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13626__A1 (.I(_03316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13626__A2 (.I(_04163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13626__A3 (.I(_05208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13627__A3 (.I(_05487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13628__A1 (.I(_05630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13628__A2 (.I(_05631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13628__A3 (.I(_05632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13629__A1 (.I(_05629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13633__A1 (.I(_05604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13638__A1 (.I(_05553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13639__A3 (.I(_05643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13640__B (.I(_05643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13643__A1 (.I(_05647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13644__A1 (.I(_03251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13644__A2 (.I(_03376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13647__A1 (.I(_05547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13648__I (.I(_01822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13649__A1 (.I(_03251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13650__A1 (.I(_05527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13650__A2 (.I(_05530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13651__A1 (.I(_05553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13652__A1 (.I(_05553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13654__C (.I(_05643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13655__A1 (.I(_05568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13659__I (.I(_05570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13660__A1 (.I(_04645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13661__A1 (.I(_04562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13663__A1 (.I(_05584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13666__A1 (.I(_04500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13668__A1 (.I(_04578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13668__A2 (.I(_05671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13670__A1 (.I(_04211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13670__A2 (.I(_05671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13676__A1 (.I(_05604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13678__A1 (.I(_05594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13679__A1 (.I(_05591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13680__A1 (.I(_04512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13680__A2 (.I(_04447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13683__I (.I(_05588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13684__A1 (.I(_04176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13685__A2 (.I(_05260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13686__S (.I(_05179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13687__A1 (.I(_04400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13687__A2 (.I(_05690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13690__A1 (.I(_05596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13690__A2 (.I(_05597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13691__A1 (.I(_05596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13691__A2 (.I(_05597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13694__A1 (.I(_04694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13694__A2 (.I(_05075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13695__A1 (.I(_04222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13697__A3 (.I(_05700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13698__A1 (.I(_05686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13705__A2 (.I(_05621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13706__A2 (.I(_05621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13708__A2 (.I(_04924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13709__A1 (.I(_04452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13709__A2 (.I(_04713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13711__A3 (.I(_05714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13714__A1 (.I(_05629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13716__A1 (.I(_04802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13716__A2 (.I(_04753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13717__I (.I(_04825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13718__A1 (.I(_03383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13718__A3 (.I(_05721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13719__A1 (.I(_03398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13719__A2 (.I(_04403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13719__A3 (.I(_04805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13720__A2 (.I(_05723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13722__A1 (.I(_05631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13722__A2 (.I(_05632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13723__A1 (.I(_05631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13723__A2 (.I(_05632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13724__A1 (.I(_05630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13725__A1 (.I(_04274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13726__A1 (.I(_03333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13728__I (.I(_05731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13729__A1 (.I(_03350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13729__A2 (.I(_04192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13730__A1 (.I(_05730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13743__A1 (.I(_05743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13743__A2 (.I(_05746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13744__A1 (.I(_05657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13745__A2 (.I(_05657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13750__A2 (.I(_03346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13756__A1 (.I(_05547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13763__I (.I(_05671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13764__A1 (.I(_04667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13765__A1 (.I(_05563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13767__A1 (.I(_05686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13770__A1 (.I(_04630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13773__A1 (.I(_04597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13775__A1 (.I(_04764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13783__I (.I(_05700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13787__A1 (.I(_04966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13787__A2 (.I(_04447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13790__I (.I(_05690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13791__A1 (.I(_04525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13792__A1 (.I(_04200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13793__S (.I(_03187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13794__A1 (.I(_04487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13794__A2 (.I(_05796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13796__A1 (.I(_05794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13797__I (.I(_04471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13798__A1 (.I(_05512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13799__A1 (.I(_04694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13801__A1 (.I(_04705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13801__A2 (.I(_05260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13802__A1 (.I(_04728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13802__A2 (.I(_05078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13803__A1 (.I(_04221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13803__A2 (.I(_05187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13805__A1 (.I(_05803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13805__A2 (.I(_05807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13807__A1 (.I(_05792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13811__A2 (.I(_05714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13812__A2 (.I(_05714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13814__A2 (.I(_05723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13815__A2 (.I(_05723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13817__A1 (.I(_05158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13817__A2 (.I(_05074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13818__A1 (.I(_04451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13818__A2 (.I(_05516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13819__A1 (.I(_04893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13825__I (.I(_05469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13827__A1 (.I(_04864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13827__A2 (.I(_05721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13828__A1 (.I(_04753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13830__A1 (.I(_05730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13832__A1 (.I(_04397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13832__A2 (.I(_04818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13833__A3 (.I(_05145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13834__A3 (.I(_05731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13841__A2 (.I(_05813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13841__A3 (.I(_05843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13846__A1 (.I(_05846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13846__A2 (.I(_05848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13847__A1 (.I(_05743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13847__A2 (.I(_05746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13849__A1 (.I(_05849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13850__I (.I(_03376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13852__A1 (.I(_03284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13853__A1 (.I(_05852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13860__A1 (.I(_05547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13861__A1 (.I(_03284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13862__A1 (.I(_05852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13866__A1 (.I(_05852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13868__A2 (.I(_05643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13869__A3 (.I(_05849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13870__A2 (.I(_05657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13870__A3 (.I(_05849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13871__A1 (.I(_05743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13871__A2 (.I(_05746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13872__A1 (.I(_05846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13872__A2 (.I(_05848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13873__A1 (.I(_05846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13873__A2 (.I(_05848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13882__A1 (.I(_04667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13883__A1 (.I(_05440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13885__A1 (.I(_05792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13888__A1 (.I(_04561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13890__I (.I(_05891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13891__A1 (.I(_04597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13893__A1 (.I(_04642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13899__A1 (.I(_05813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13899__A2 (.I(_05843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13900__A1 (.I(_05813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13900__A2 (.I(_05843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13907__I (.I(_05229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13908__A1 (.I(_04406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13908__A2 (.I(_05909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13908__B2 (.I(_04929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13909__A1 (.I(_04406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13909__A2 (.I(_04929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13911__A1 (.I(_04324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13911__A2 (.I(_05078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13912__A1 (.I(_04451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13913__A2 (.I(_04927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13921__A2 (.I(_05208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13922__A2 (.I(_05731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13923__A2 (.I(_04818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13927__A2 (.I(_05229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13934__A1 (.I(_05803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13934__A2 (.I(_05807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13936__A1 (.I(_04446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13936__A2 (.I(_04766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13939__A1 (.I(_04176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13939__A2 (.I(_05796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13940__A2 (.I(_05504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13941__I1 (.I(\filters.band[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13941__S (.I(_05179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13942__A1 (.I(_04186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13942__A2 (.I(_05943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13946__A1 (.I(_04238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13946__B2 (.I(_04847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13947__A1 (.I(_04238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13947__A2 (.I(_04847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13949__A1 (.I(_04229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13950__A1 (.I(_04254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13950__A2 (.I(_05185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13951__A1 (.I(_04392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13953__A1 (.I(_05950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13953__A2 (.I(_05954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13955__A1 (.I(_05940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13957__A1 (.I(_05905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13957__A2 (.I(_05935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13966__A1 (.I(_05877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13966__A2 (.I(_05967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13967__I (.I(\filters.low[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13968__A1 (.I(_05969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13969__A1 (.I(_03299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13970__A1 (.I(_05968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13974__I (.I(_05543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13980__A1 (.I(_05560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13981__I (.I(_04631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13982__A1 (.I(_05982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13984__A1 (.I(_05940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13987__A1 (.I(_04630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13988__I (.I(_05796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13990__A1 (.I(_04616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13990__A2 (.I(_05990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13992__A1 (.I(_04498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13992__A2 (.I(_05990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13997__A1 (.I(_05905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13997__A2 (.I(_05935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13998__A1 (.I(_05905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13998__A2 (.I(_05935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14000__A1 (.I(_05950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14000__A2 (.I(_05954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14004__I (.I(_05943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14005__A1 (.I(_04529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14006__A1 (.I(_04742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14006__A2 (.I(_05588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14007__I0 (.I(\filters.high[25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14007__I1 (.I(\filters.band[25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14007__S (.I(_03187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14008__A1 (.I(_04487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14008__A2 (.I(_06008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14011__A1 (.I(_05512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14012__A1 (.I(_04694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14014__A1 (.I(_04728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14015__A1 (.I(_04259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14017__A1 (.I(_06015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14017__A2 (.I(_06016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14018__A1 (.I(_06014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14020__A1 (.I(_06004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14027__A1 (.I(_04397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14027__B1 (.I(_06027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14028__A2 (.I(_04397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14028__A4 (.I(_06027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14030__A2 (.I(_04341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14031__A2 (.I(_04403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14033__A1 (.I(_04750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14033__A2 (.I(_04884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14035__A1 (.I(_06030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14037__A1 (.I(_05469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14037__A2 (.I(_04825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14038__A1 (.I(_05516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14041__A2 (.I(_06041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14045__A1 (.I(_04929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14046__A3 (.I(_05721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14048__A1 (.I(_04377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14048__A2 (.I(_05074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14049__A1 (.I(_04372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14049__A2 (.I(_05078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14055__A1 (.I(_06024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14055__A2 (.I(_06055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14063__A1 (.I(_05877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14063__A2 (.I(_05967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14063__B (.I(net46));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14064__A1 (.I(_06062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14067__A1 (.I(_03310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14067__A2 (.I(_03377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14068__A1 (.I(_03314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14068__A2 (.I(_06067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14069__A1 (.I(_06065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14070__A1 (.I(_06065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14072__I (.I(_03472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14073__A1 (.I(_03299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14073__A2 (.I(_06073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14073__B (.I(_05968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14079__A1 (.I(_03314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14080__I (.I(_05544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14086__I (.I(_05990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14087__A1 (.I(_04645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14088__A1 (.I(_05440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14091__A1 (.I(_06004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14092__A1 (.I(_04561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14094__A1 (.I(_05446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14097__A1 (.I(_04416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14102__A1 (.I(_06024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14102__A2 (.I(_06055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14104__A2 (.I(_06041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14106__A1 (.I(_06030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14110__A3 (.I(_05106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14111__A1 (.I(_03413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14111__A2 (.I(_04488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14113__A1 (.I(_04711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14116__A1 (.I(_04740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14116__A2 (.I(_04781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14117__A1 (.I(_04803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14119__A2 (.I(_04927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14129__A1 (.I(_04376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14129__A2 (.I(_05077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14130__A1 (.I(_04371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14130__A2 (.I(_05185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14131__A1 (.I(_04367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14136__A1 (.I(_06105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14136__A2 (.I(_06135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14137__A1 (.I(_06014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14143__A1 (.I(_04529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14143__A2 (.I(_06008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14144__A1 (.I(_04742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14144__A2 (.I(_05690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14145__A1 (.I(\filters.band[26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14145__A2 (.I(_04186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14148__A1 (.I(_06015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14148__A2 (.I(_06016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14149__A1 (.I(_06015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14149__A2 (.I(_06016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14151__A1 (.I(_05069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14151__A2 (.I(_05350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14152__A1 (.I(_04258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14152__A2 (.I(_05504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14154__A2 (.I(_05588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14156__A2 (.I(_06155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14158__A1 (.I(_06142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14169__A1 (.I(_05967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14169__A2 (.I(_06062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14174__I (.I(_06173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14175__A1 (.I(_05877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14176__A1 (.I(_06168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14178__A1 (.I(_03329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14179__A1 (.I(_03330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14179__A2 (.I(_06177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14180__A2 (.I(_06179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14186__I (.I(_01821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14187__I (.I(_06186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14188__A1 (.I(_03330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14194__A1 (.I(_06105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14194__A2 (.I(_06135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14206__A1 (.I(_04750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14207__A1 (.I(_04737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14207__A2 (.I(_05731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14212__A2 (.I(_05049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14213__A2 (.I(_05075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14214__A1 (.I(_04896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14214__A2 (.I(_05181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14215__A1 (.I(_06211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14223__A1 (.I(_04326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14224__A1 (.I(_04452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14225__A1 (.I(_04893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14231__A1 (.I(_06197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14231__A2 (.I(_06229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14232__A2 (.I(_06155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14238__A1 (.I(\filters.band[26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14238__A2 (.I(_04596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14239__A1 (.I(_04504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14240__A1 (.I(\filters.band[27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14244__A1 (.I(_04699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14245__A1 (.I(_04697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14247__A1 (.I(_04231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14247__A2 (.I(_05891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14251__A1 (.I(_06236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14251__A2 (.I(_06249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14255__I (.I(_05560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14257__A1 (.I(_05982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14259__A1 (.I(_06142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14262__I (.I(_06008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14263__A1 (.I(_04616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14263__A2 (.I(_06261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14265__A1 (.I(_04644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14265__A2 (.I(_06261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14267__A1 (.I(_05440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14276__A2 (.I(_06192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14279__A1 (.I(_06275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14279__A2 (.I(_06277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14280__I (.I(_06168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14283__B (.I(_06281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14285__A1 (.I(_03345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14286__A1 (.I(_03347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14286__A2 (.I(_06177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14287__A2 (.I(_06285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14289__A2 (.I(_06179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14290__A2 (.I(_06179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14294__A1 (.I(_03347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14297__A2 (.I(_06285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14298__A2 (.I(_06179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14298__B2 (.I(_06285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14301__A1 (.I(_06168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14303__A1 (.I(_06275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14303__A2 (.I(_06277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14304__A1 (.I(_06281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14304__B2 (.I(_06173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14305__A1 (.I(_06275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14305__A2 (.I(_06277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14306__A1 (.I(_05877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14311__A1 (.I(_06197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14311__A2 (.I(_06229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14322__A1 (.I(_05469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14322__A2 (.I(_06027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14323__A1 (.I(_04858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14323__A2 (.I(_05487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14325__A2 (.I(_04924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14328__A1 (.I(_05909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14328__A2 (.I(_05092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14329__A1 (.I(_04806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14330__A1 (.I(_04446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14334__I (.I(_04355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14335__A2 (.I(_05570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14337__A1 (.I(_06211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14338__A1 (.I(_06211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14340__A1 (.I(_04326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14341__A1 (.I(_04378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14342__A1 (.I(_04318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14345__A1 (.I(_06337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14349__A1 (.I(_06314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14349__A2 (.I(_06346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14356__A1 (.I(\filters.band[27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14356__A2 (.I(_04578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14359__A2 (.I(_04617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14362__A2 (.I(_05891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14365__A1 (.I(_05509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14366__A1 (.I(_04222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14373__A2 (.I(_06370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14376__A1 (.I(_06236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14376__A2 (.I(_06249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14382__I (.I(\filters.band[26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14383__A2 (.I(_04632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14385__I (.I(_06261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14386__A1 (.I(_05563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14389__A1 (.I(_06373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14391__A1 (.I(_06308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14392__A1 (.I(_06305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14393__A1 (.I(_06192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14394__A1 (.I(_06192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14397__A2 (.I(_06394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14400__A1 (.I(_03360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14400__A2 (.I(_03221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14401__A1 (.I(_03361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14401__A2 (.I(_06397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14402__A2 (.I(_06399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14403__A1 (.I(_06298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14405__A1 (.I(_03361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14406__I (.I(_05543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14408__A1 (.I(_06373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14413__A1 (.I(_06314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14413__A2 (.I(_06346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14414__A2 (.I(_06370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14424__A2 (.I(_06027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14426__A2 (.I(_05075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14428__A1 (.I(_06420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14429__A1 (.I(_05721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14430__A1 (.I(_04805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14430__A2 (.I(_05187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14432__A1 (.I(_04802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14435__A1 (.I(_06417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14435__A2 (.I(_06431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14437__A2 (.I(_05671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14442__A1 (.I(_04355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14443__A1 (.I(_04453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14444__A1 (.I(_04318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14456__A1 (.I(_06337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14457__A2 (.I(_05446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14458__A2 (.I(_06261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14460__A1 (.I(_06456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14460__A2 (.I(_04617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14462__A1 (.I(_04576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14462__A2 (.I(_05990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14465__A1 (.I(_05509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14466__A1 (.I(_05510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14477__A1 (.I(_06472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14478__A1 (.I(_05982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14483__A2 (.I(_05563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14487__I (.I(\filters.band[27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14488__A2 (.I(_05560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14494__A1 (.I(_06308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14495__A1 (.I(_06305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14498__A2 (.I(_06394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14503__A1 (.I(_03374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14503__A2 (.I(_06177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14504__A1 (.I(_03380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14504__A2 (.I(_03378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14505__A2 (.I(_06501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14506__A2 (.I(_06399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14507__A1 (.I(_06298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14510__A1 (.I(_06403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14511__A1 (.I(_03380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14512__I (.I(_05544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14525__A1 (.I(_06520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14531__A2 (.I(_04631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14535__A2 (.I(_04667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14547__A2 (.I(_05446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14549__A1 (.I(\filters.band[30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14549__A2 (.I(_04506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14556__A2 (.I(_06008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14557__A1 (.I(_05512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14557__A2 (.I(_05796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14558__A1 (.I(_05510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14565__A1 (.I(_06417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14565__A2 (.I(_06431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14568__A1 (.I(_04355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14570__A1 (.I(_04446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14572__A1 (.I(_04326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14572__A2 (.I(_05891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14573__A1 (.I(_04452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14574__A1 (.I(_04893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14579__A1 (.I(_06420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14581__A1 (.I(_04802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14582__A1 (.I(_05909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14583__A1 (.I(_04806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14589__A1 (.I(_04924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14589__A2 (.I(_05626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14590__A1 (.I(_05624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14604__A2 (.I(_03377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14605__A1 (.I(_03396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14605__A2 (.I(_06067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14606__A1 (.I(_06599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14606__A2 (.I(_06601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14608__A2 (.I(_06501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14609__A2 (.I(_06501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14611__A1 (.I(_06298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14613__A1 (.I(_06403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14614__I (.I(_06186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14615__A1 (.I(_03396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14620__A1 (.I(_06614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14623__A1 (.I(_04222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14624__A1 (.I(_06520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14624__A2 (.I(_04601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14628__A1 (.I(_05909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14633__A1 (.I(_04318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14634__A1 (.I(_04447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14635__A1 (.I(_05624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14635__A2 (.I(_05281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14641__A3 (.I(_06635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14645__A1 (.I(_06472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14645__A2 (.I(_04576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14646__A1 (.I(_04576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14648__A1 (.I(_05509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14652__A1 (.I(\filters.band[31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14658__A1 (.I(_06614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14658__A2 (.I(_05982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14668__A1 (.I(_06456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14673__A1 (.I(_04806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14675__A1 (.I(_05268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14675__A2 (.I(_05626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14680__A1 (.I(\filters.band[30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14682__A1 (.I(_04453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14685__A1 (.I(_06675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14689__A2 (.I(_06682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14694__I (.I(_06688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14695__A1 (.I(_03411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14695__A2 (.I(_03221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14696__A1 (.I(_03412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14696__A2 (.I(_03378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14697__A1 (.I(_06689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14697__A2 (.I(_06691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14698__A1 (.I(_06599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14698__A2 (.I(_06601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14706__I (.I(_06688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14708__A1 (.I(_06701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14708__A2 (.I(_06691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14710__A1 (.I(_06703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14710__A2 (.I(_06691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14713__A1 (.I(_06706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14713__A2 (.I(_06691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14715__A1 (.I(_06298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14716__I (.I(_06067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14717__A1 (.I(_03422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14717__A2 (.I(_06397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14718__A2 (.I(_06710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14719__A1 (.I(_06689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14719__A2 (.I(_06712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14721__A1 (.I(\filters.band[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14722__A2 (.I(_06714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14723__I (.I(_06703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14725__I (.I(_06717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14728__A1 (.I(_06720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14728__A2 (.I(_06712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14730__A1 (.I(_06722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14730__A2 (.I(_06712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14732__A2 (.I(_06710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14734__A1 (.I(_06689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14736__A1 (.I(_06403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14738__A2 (.I(_06397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14740__A1 (.I(_06703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14740__A2 (.I(_06731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14743__A1 (.I(_06712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14743__B (.I(_06734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14746__A1 (.I(_06403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14749__A1 (.I(_03468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14749__A2 (.I(_06710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14751__A2 (.I(_06703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14752__A1 (.I(_06722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14752__A2 (.I(_06731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14756__A1 (.I(_05544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14758__I (.I(_05546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14761__A1 (.I(_06731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14761__B (.I(_06734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14763__I (.I(_06752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14765__I (.I(_03472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14766__I0 (.I(\filters.low[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14766__I1 (.I(\filters.band[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14770__I (.I(_04159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14771__I (.I(_06760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14772__I (.I(_03733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14774__A1 (.I(\filters.band[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14774__A2 (.I(_06761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14777__I (.I(_06765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14781__A1 (.I(_06769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14783__I0 (.I(\filters.low[17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14786__I (.I(_03721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14787__A2 (.I(_04160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14787__B (.I(_06775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14788__A1 (.I(_06761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14789__I (.I(_06689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14790__I1 (.I(\filters.band[18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14790__S (.I(_06073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14792__B (.I(_06765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14797__I (.I(_06760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14798__A1 (.I(\filters.band[18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14801__A1 (.I(_06706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14803__A1 (.I(_06769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14808__S (.I(_03472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14809__A1 (.I(_06701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14812__B (.I(_06734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14819__I (.I(_05546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14821__A1 (.I(_06769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14822__I1 (.I(\filters.band[21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14822__S (.I(_06073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14827__A1 (.I(\filters.band[21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14829__S (.I(_06073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14832__B (.I(_06765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14836__I (.I(_06760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14841__A2 (.I(_03473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14843__A1 (.I(_06720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14851__B (.I(_06717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14853__B2 (.I(_06752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14854__I (.I(_06701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14856__A1 (.I(\filters.band[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14860__A1 (.I(\filters.band[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14860__A2 (.I(_04160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14860__B (.I(_06775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14861__A1 (.I(_06761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14863__A1 (.I(_06722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14865__I1 (.I(\filters.band[25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14865__S (.I(_03473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14869__A1 (.I(\filters.band[25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14871__I (.I(_05546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14872__I (.I(_06706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14873__I1 (.I(_06472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14873__S (.I(_03473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14881__A1 (.I(_06472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14883__I (.I(_06706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14884__I1 (.I(_06520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14890__I (.I(_06760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14891__A1 (.I(_06520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14898__A1 (.I(_06614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14899__A2 (.I(_03476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14903__A1 (.I(_06614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14906__A1 (.I(_06456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14913__A1 (.I(_06456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14914__A1 (.I(_06889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14916__A1 (.I(\filters.band[30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14916__A2 (.I(_03476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14921__A1 (.I(_06722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14922__A1 (.I(_05547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14924__A1 (.I(\filters.band[30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14924__B (.I(_06899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14926__A1 (.I(_06720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14927__A1 (.I(_06720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14929__I1 (.I(\filters.band[31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14930__A1 (.I(_06769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14931__A1 (.I(\filters.band[31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14931__A2 (.I(_04160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14931__B (.I(_06775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14932__A1 (.I(_06761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14933__A1 (.I(_03730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14933__A2 (.I(_04170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14936__I (.I(_06909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14940__A2 (.I(_06912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14940__B (.I(_06913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14942__A1 (.I(_05534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14942__A2 (.I(_06915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14944__A2 (.I(_06910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14944__C (.I(_06917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14945__I (.I(_01932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14949__A3 (.I(\channels.sample1[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14949__A4 (.I(\channels.sample2[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14950__A2 (.I(\channels.sample1[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14950__B1 (.I(\channels.sample2[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14952__A2 (.I(\channels.sample3[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14953__A1 (.I(_05647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14955__A2 (.I(_06912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14956__A1 (.I(_05534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14956__A2 (.I(_06915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14957__A1 (.I(_06921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14958__B (.I(_06921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14959__A1 (.I(_06909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14960__A1 (.I(\filters.high[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14960__A2 (.I(_06919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14965__A1 (.I(_01773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14965__A2 (.I(\channels.sample3[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14966__A1 (.I(_05647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14968__A3 (.I(\channels.sample1[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14968__A4 (.I(\channels.sample2[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14969__A2 (.I(\channels.sample1[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14969__B1 (.I(\channels.sample2[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14971__A2 (.I(\channels.sample3[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14977__A2 (.I(_05035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14978__A2 (.I(_06949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14981__B (.I(_06952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14982__A1 (.I(\filters.high[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14982__A2 (.I(_06934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14984__I (.I(_06952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14985__A1 (.I(\filters.high[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14985__A2 (.I(_06955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14986__A2 (.I(_06949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14991__A1 (.I(\filters.filt_2 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14991__A2 (.I(\filters.filt_1 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14991__A3 (.I(\channels.sample1[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14991__A4 (.I(\channels.sample2[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14992__A1 (.I(\filters.filt_1 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14992__A2 (.I(\channels.sample1[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14992__B1 (.I(\channels.sample2[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14992__B2 (.I(\filters.filt_2 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14994__A1 (.I(\filters.filt_3 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14994__A2 (.I(\channels.sample3[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14999__A2 (.I(_05035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15001__A2 (.I(_05035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15005__B (.I(_06952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15007__I (.I(_03940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15008__I (.I(_06978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15009__B (.I(_06979_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15010__A2 (.I(_06955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15011__A1 (.I(_04158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15011__A2 (.I(_04776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15017__A1 (.I(\filters.filt_2 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15017__A2 (.I(\filters.filt_1 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15017__A3 (.I(\channels.sample1[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15017__A4 (.I(\channels.sample2[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15018__A2 (.I(\channels.sample1[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15018__B1 (.I(\channels.sample2[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15020__A2 (.I(\channels.sample3[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15027__A1 (.I(\filters.low[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15027__A3 (.I(_06996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15035__A1 (.I(_06983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15036__B (.I(_06979_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15039__A1 (.I(_05969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15040__A1 (.I(_05969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15041__A2 (.I(_06996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15042__B (.I(_04993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15049__A2 (.I(\channels.sample3[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15050__A2 (.I(\channels.sample2[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15051__A2 (.I(\channels.sample1[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15056__A1 (.I(_04992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15062__B (.I(_07030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15065__A1 (.I(\filters.high[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15065__A2 (.I(_07033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15065__B (.I(_06899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15066__A1 (.I(_07032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15067__I (.I(_07030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15077__A2 (.I(\channels.sample2[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15078__A2 (.I(\channels.sample1[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15088__A1 (.I(_04992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15089__A1 (.I(_03310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15095__A1 (.I(\filters.high[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15095__A2 (.I(_07062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15095__B (.I(_06775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15096__A2 (.I(_07061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15097__I (.I(_06913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15098__A1 (.I(_05417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15098__A2 (.I(_05420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15103__A2 (.I(_01927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15106__A2 (.I(\channels.sample3[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15107__A2 (.I(\channels.sample2[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15108__A2 (.I(\channels.sample1[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15113__A1 (.I(_03329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15120__B (.I(_07086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15122__I (.I(_06186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15141__A2 (.I(\channels.sample2[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15142__A2 (.I(\channels.sample1[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15149__A1 (.I(_03345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15154__A1 (.I(_06913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15154__A2 (.I(_07119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15156__A1 (.I(_05379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15156__A2 (.I(_05403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15161__A2 (.I(_01977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15164__A2 (.I(\channels.sample3[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15165__A2 (.I(\channels.sample2[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15166__A2 (.I(\channels.sample1[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15169__A2 (.I(_07133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15170__A2 (.I(_07122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15172__A1 (.I(_03360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15177__B (.I(_07086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15194__A2 (.I(\channels.sample2[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15195__A2 (.I(\channels.sample1[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15199__A3 (.I(_07162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15201__A2 (.I(_07122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15203__A1 (.I(_03374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15203__A2 (.I(_07133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15205__A2 (.I(_07168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15206__A1 (.I(_07146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15206__A2 (.I(_07149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15207__A2 (.I(_07146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15207__A3 (.I(_07149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15208__A1 (.I(_06909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15209__A1 (.I(\filters.high[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15209__A2 (.I(_06934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15211__A1 (.I(_03394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15211__A2 (.I(_07162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15212__A1 (.I(_03394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15212__A2 (.I(_07162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15217__A2 (.I(_02029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15220__A2 (.I(\channels.sample3[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15221__A1 (.I(_01762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15221__A2 (.I(\channels.sample2[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15222__A1 (.I(_01748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15222__A2 (.I(\channels.sample1[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15225__A2 (.I(_07187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15226__A1 (.I(_03411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15226__A2 (.I(_07187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15230__A2 (.I(_07168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15231__B (.I(_07086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15233__A1 (.I(_03410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15235__A1 (.I(_07146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15235__A2 (.I(_07149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15236__A2 (.I(_07168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15249__A2 (.I(\channels.sample3[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15250__A2 (.I(\channels.sample2[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15251__A2 (.I(\channels.sample1[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15255__A2 (.I(_07216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15256__A1 (.I(_03422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15256__A2 (.I(_07216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15261__I (.I(_03721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15262__A1 (.I(\filters.high[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15262__A2 (.I(_07062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15265__A2 (.I(_02056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15270__A1 (.I(_07227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15270__A2 (.I(_07230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15273__A1 (.I(_05849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15273__A3 (.I(_07233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15280__B (.I(_07240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15282__A2 (.I(_07033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15282__B (.I(_06899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15284__A1 (.I(_07227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15284__A2 (.I(_07230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15286__A1 (.I(_05968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15289__A1 (.I(_05852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15289__A2 (.I(_07233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15299__A2 (.I(_06955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15301__A2 (.I(_06065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15302__A1 (.I(_05968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15308__B (.I(_07086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15310__I (.I(_06186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15311__A2 (.I(_06910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15311__C (.I(_07269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15320__A1 (.I(_03468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15320__A2 (.I(_06065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15321__A1 (.I(\filters.low[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15323__A1 (.I(_07277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15324__A2 (.I(_07062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15326__A1 (.I(\filters.low[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15327__A1 (.I(\filters.low[17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15329__A1 (.I(_07277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15331__A1 (.I(_06919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15332__A2 (.I(_07033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15332__B (.I(_06899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15334__A2 (.I(_06955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15335__A1 (.I(\filters.low[17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15339__I (.I(\filters.low[17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15340__A1 (.I(_07295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15344__A1 (.I(_07277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15346__A1 (.I(_06983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15347__B (.I(_06979_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15351__A1 (.I(_07295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15352__A1 (.I(_07295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15358__I (.I(_07030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15360__A2 (.I(_06599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15367__B2 (.I(_07277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15368__A2 (.I(_07321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15372__A2 (.I(_07321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15375__A2 (.I(_06599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15377__B (.I(_07240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15379__I (.I(_03733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15380__I (.I(_07332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15381__A2 (.I(_07033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15381__B (.I(_07333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15383__A2 (.I(_06919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15389__A1 (.I(_07321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15395__A1 (.I(_07062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15396__B (.I(_06979_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15401__A2 (.I(_06701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15405__I (.I(_07355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15406__B (.I(_07356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15412__B2 (.I(_07321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15418__B (.I(_07356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15420__I (.I(\filters.high[25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15429__A1 (.I(_07373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15432__A1 (.I(_06934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15433__A2 (.I(_06910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15433__C (.I(_06917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15434__I (.I(_01932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15437__A2 (.I(_06765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15441__A1 (.I(_07373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15445__A1 (.I(_06909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15446__A2 (.I(_06934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15450__A2 (.I(_06734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15452__A1 (.I(_07373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15454__B (.I(_07240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15456__A2 (.I(_06983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15456__B (.I(_07333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15464__A2 (.I(_06717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15468__A2 (.I(_07030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15468__B (.I(_07356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15469__A2 (.I(_07413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15472__A2 (.I(_06717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15476__B (.I(_07240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15478__A2 (.I(_06983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15478__B (.I(_07333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15480__A2 (.I(_06919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15489__B (.I(_06952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15491__I (.I(_06978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15499__B (.I(_06913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15500__A2 (.I(_06910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15500__C (.I(_06917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15501__I (.I(_03202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15502__A1 (.I(\filters.mode_vol[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15502__A2 (.I(_01773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15502__C (.I(_03215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15503__A1 (.I(_01748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15503__B1 (.I(_03476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15503__B2 (.I(_01762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15504__C (.I(_03729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15505__I (.I(_07446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15507__A1 (.I(_03194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15507__A2 (.I(_04189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15507__B (.I(_07446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15510__A1 (.I(_03202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15510__A2 (.I(_03204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15510__A3 (.I(_03215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15512__A1 (.I(\channels.sample3[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15513__A1 (.I(_03263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15514__A1 (.I(\channels.sample2[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15515__A1 (.I(\channels.sample1[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15517__A2 (.I(_07458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15520__I (.I(_07446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15521__A2 (.I(_07458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15523__A1 (.I(\channels.sample3[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15525__A1 (.I(\channels.sample2[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15526__A1 (.I(\channels.sample1[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15528__A2 (.I(_07468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15532__A2 (.I(_07468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15534__A1 (.I(\channels.sample3[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15536__A1 (.I(\channels.sample2[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15536__A2 (.I(_03346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15537__A1 (.I(\channels.sample1[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15539__A2 (.I(_07478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15545__I (.I(_07446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15546__A1 (.I(\filters.sample_buff[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15548__A2 (.I(_07478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15550__A1 (.I(\channels.sample3[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15551__C (.I(_03376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15552__A1 (.I(\channels.sample2[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15553__A1 (.I(\channels.sample1[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15555__A1 (.I(\filters.sample_buff[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15555__A2 (.I(_07493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15560__I (.I(_01932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15561__A1 (.I(\filters.sample_buff[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15561__A2 (.I(_07493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15562__A1 (.I(\channels.sample3[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15564__A1 (.I(\channels.sample2[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15564__A2 (.I(_03377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15565__A1 (.I(\channels.sample1[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15567__A1 (.I(\filters.sample_buff[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15567__A2 (.I(_07504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15572__A1 (.I(\filters.sample_buff[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15575__A1 (.I(\filters.sample_buff[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15575__A2 (.I(_07504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15577__A1 (.I(_01927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15578__C (.I(_06067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15579__A1 (.I(\channels.sample2[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15579__A2 (.I(_03378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15580__A1 (.I(\channels.sample1[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15582__A2 (.I(_07518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15588__A2 (.I(_07518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15589__A1 (.I(\channels.sample3[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15590__C (.I(_06177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15591__A1 (.I(\channels.sample2[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15591__A2 (.I(_06397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15592__A1 (.I(\channels.sample1[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15594__A2 (.I(_07529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15602__A2 (.I(_07529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15604__A1 (.I(_01977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15605__C (.I(_06710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15606__A1 (.I(\channels.sample2[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15606__A2 (.I(_03395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15607__A1 (.I(\channels.sample1[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15609__A2 (.I(_07543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15614__A2 (.I(_07543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15616__A1 (.I(\channels.sample3[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15617__C (.I(_03395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15618__A1 (.I(\channels.sample2[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15619__A1 (.I(\channels.sample1[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15621__A2 (.I(_07554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15629__A2 (.I(_07554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15631__A1 (.I(_02029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15633__A1 (.I(\channels.sample2[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15634__A1 (.I(\channels.sample1[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15636__A2 (.I(_07568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15640__I (.I(_06978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15641__B (.I(_07573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15642__A2 (.I(_07568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15643__A1 (.I(\channels.sample3[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15645__A1 (.I(\channels.sample2[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15646__A1 (.I(\channels.sample1[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15648__A1 (.I(\filters.sample_buff[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15648__A2 (.I(_07579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15653__A1 (.I(\filters.sample_buff[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15655__A1 (.I(\filters.sample_buff[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15656__A1 (.I(\filters.sample_buff[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15656__A2 (.I(_07579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15657__A1 (.I(_02056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15659__A1 (.I(\channels.sample2[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15660__A1 (.I(\channels.sample1[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15662__A1 (.I(\filters.sample_buff[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15662__A2 (.I(_07592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15666__B (.I(_07573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15667__I (.I(_03940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15669__A1 (.I(\filters.sample_buff[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15669__A2 (.I(_07592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15671__A1 (.I(_03239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15673__A1 (.I(\filters.sample_buff[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15674__B (.I(\filters.sample_buff[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15677__A1 (.I(\filters.sample_buff[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15678__A1 (.I(_07598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15679__A1 (.I(\filters.sample_buff[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15682__A1 (.I(\filters.sample_buff[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15686__B (.I(_07573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15688__A1 (.I(\filters.sample_buff[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15695__C (.I(_07269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15706__A2 (.I(_03729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15709__I (.I(_07630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15710__I (.I(_07631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15711__I (.I(_07630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15712__A1 (.I(_05534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15712__B (.I(_07356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15713__A2 (.I(_07632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15714__A2 (.I(_03730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15714__A3 (.I(_03205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15715__I (.I(_07635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15716__I (.I(_07636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15719__I (.I(_07639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15720__A1 (.I(_05647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15720__A2 (.I(_07640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15720__B (.I(_07333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15723__I (.I(_07639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15724__I (.I(_07332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15730__I (.I(_07355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15731__A1 (.I(_05969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15731__B (.I(_07648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15732__A2 (.I(_07632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15734__A1 (.I(_03310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15735__A1 (.I(_07650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15736__I (.I(_07636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15738__A1 (.I(_03329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15739__A1 (.I(_07653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15741__I (.I(_07639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15742__I (.I(_07332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15743__A1 (.I(_03345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15746__A1 (.I(_03360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15747__A1 (.I(_07659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15749__A1 (.I(_03374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15751__I (.I(_07635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15752__I (.I(_07663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15754__A1 (.I(_03394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15755__A1 (.I(_07665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15756__A1 (.I(_03411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15756__B (.I(_07648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15757__A2 (.I(_07632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15758__A1 (.I(_03422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15758__B (.I(_07648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15759__A1 (.I(_06714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15759__A2 (.I(_07632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15761__I (.I(_07639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15762__I (.I(_07332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15763__A2 (.I(_07670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15763__B (.I(_07671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15766__A2 (.I(_07670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15766__B (.I(_07671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15769__A1 (.I(_03468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15769__A2 (.I(_07670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15769__B (.I(_07671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15771__I (.I(_07663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15773__A1 (.I(\filters.low[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15773__A2 (.I(_07670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15773__B (.I(_07671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15775__A1 (.I(_07295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15775__A2 (.I(_07631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15775__B (.I(_07648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15776__A2 (.I(_07640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15778__I (.I(_07630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15779__I (.I(_03733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15780__I (.I(_07683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15781__A2 (.I(_07682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15781__B (.I(_07684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15784__A2 (.I(_07682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15784__B (.I(_07684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15787__A2 (.I(_07682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15787__B (.I(_07684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15789__I (.I(_07663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15791__A2 (.I(_07682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15791__B (.I(_07684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15794__I (.I(_07630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15795__I (.I(_07683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15798__I (.I(_07636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15799__I (.I(_07663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15801__A2 (.I(_07697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15801__C (.I(_07269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15802__I (.I(_07355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15803__A2 (.I(_07631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15803__B (.I(_07700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15804__A2 (.I(_07640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15806__A1 (.I(_07373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15815__A2 (.I(_07697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15815__C (.I(_07269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15818__A2 (.I(_07697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15818__C (.I(_07710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15819__A2 (.I(_07636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15820__A2 (.I(_07697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15820__C (.I(_07710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15821__A2 (.I(_07631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15821__B (.I(_07700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15822__A2 (.I(_07640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15823__A1 (.I(_03735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15824__A1 (.I(_04189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15824__A2 (.I(_04158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15825__A3 (.I(_03731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15826__A1 (.I(_03735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15827__A1 (.I(_03194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15829__A1 (.I(_07598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15835__I (.I(_07721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15836__A2 (.I(_04776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15836__A3 (.I(_07722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15837__B (.I(_07573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15841__A2 (.I(_07726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15844__A1 (.I(_04776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15844__A2 (.I(_07721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15846__A2 (.I(_07728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15847__A1 (.I(_07598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15851__A1 (.I(_07721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15852__A1 (.I(_03735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15856__I (.I(_01822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15857__B (.I(_07740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15859__I (.I(_07741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15860__I (.I(_07742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15862__A1 (.I(_04170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15862__C (.I(_07710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15883__I (.I(\tt_um_rejunity_sn76489.chan[1].attenuation.in ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15886__A1 (.I(\tt_um_rejunity_sn76489.chan[1].attenuation.control[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15888__A1 (.I(\tt_um_rejunity_sn76489.chan[1].attenuation.control[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15890__A1 (.I(\tt_um_rejunity_sn76489.chan[1].attenuation.control[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15893__A2 (.I(\tt_um_rejunity_sn76489.chan[1].attenuation.in ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15896__A1 (.I(\tt_um_rejunity_sn76489.chan[1].attenuation.control[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15925__I (.I(_07806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15952__I (.I(_07726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15955__A2 (.I(_07728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15956__A1 (.I(_07598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15957__I (.I(_07722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15976__A1 (.I(\tt_um_rejunity_sn76489.chan[1].attenuation.control[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15990__I (.I(_02101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15992__A1 (.I(_07838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16035__A1 (.I(_07880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16035__A3 (.I(_07914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16043__A1 (.I(_07838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16055__A1 (.I(\tt_um_rejunity_sn76489.chan[1].attenuation.control[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16064__A1 (.I(_07929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16064__A3 (.I(_07942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16065__A2 (.I(_07914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16066__A2 (.I(_07914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16067__A1 (.I(_07880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16070__B (.I(_07721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16071__A2 (.I(_07726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16073__A2 (.I(_07924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16074__A1 (.I(_07923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16091__A1 (.I(_07956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16092__A2 (.I(_07942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16093__A2 (.I(_07942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16094__A1 (.I(_07929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16097__A1 (.I(_07838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16101__I (.I(_07956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16222__A1 (.I(_07726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16225__I (.I(_07683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16226__A2 (.I(_07924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16226__B (.I(_08098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16235__B (.I(_07741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16238__B (.I(_08098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16241__A2 (.I(_07722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16241__B1 (.I(_08111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16242__B (.I(_07700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16243__A1 (.I(_07924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16244__A1 (.I(\filters.sample_buff[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16244__A2 (.I(_07722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16244__B1 (.I(_07728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16245__A1 (.I(_07923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16246__I (.I(_07741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16249__A1 (.I(\filters.sample_buff[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16249__C2 (.I(_07728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16250__A1 (.I(_07923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16253__A1 (.I(_07923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16260__I (.I(_07741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16268__A1 (.I(\filters.sample_buff[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16270__A1 (.I(\filters.sample_buff[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16272__A1 (.I(\filters.sample_buff[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16272__A2 (.I(_07742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16274__A1 (.I(\filters.sample_buff[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16274__A2 (.I(_07742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16276__I (.I(_03940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16278__A2 (.I(_07742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16279__A1 (.I(_08136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16280__A1 (.I(net20));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16282__B (.I(_07740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16283__A1 (.I(net19));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16285__B (.I(_07740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16286__A1 (.I(_02103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16286__A2 (.I(_07838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16288__A1 (.I(_02354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16319__A1 (.I(_02363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16321__A1 (.I(_02363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16321__A2 (.I(_03936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16321__B (.I(_01821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16334__A1 (.I(_03964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16336__A1 (.I(_03974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16338__A1 (.I(_03978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16341__B1 (.I(_01258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16343__B1 (.I(_01258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16345__A2 (.I(_01317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16345__B1 (.I(_01258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16347__A2 (.I(_01317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16347__B1 (.I(_01334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16349__A2 (.I(_01317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16349__B1 (.I(_01334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16351__A1 (.I(_02356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16353__A1 (.I(_02356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16353__A2 (.I(_03936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16353__B (.I(_01821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16355__A1 (.I(\channels.ch3_env[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16357__A1 (.I(\channels.ch3_env[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16359__A1 (.I(\channels.ch3_env[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16361__A1 (.I(\channels.ch3_env[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16365__A1 (.I(\channels.ch3_env[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16366__A1 (.I(_03964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16367__A1 (.I(\channels.ch3_env[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16368__A1 (.I(_03974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16369__A1 (.I(\channels.ch3_env[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16370__A1 (.I(_03978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16371__A1 (.I(\channels.ch3_env[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16377__A2 (.I(_01042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16378__I (.I(_08194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16399__I (.I(_08194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16414__I (.I(_08194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16437__A2 (.I(_08238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16438__A1 (.I(_08136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16442__I (.I(_08242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16444__A2 (.I(_08244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16446__A1 (.I(_04101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16448__B (.I(_08098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16451__B (.I(_08098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16454__I (.I(_07683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16455__B (.I(_08252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16457__B (.I(_07700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16461__A1 (.I(_08136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16462__A1 (.I(_08136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16462__A2 (.I(_07924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16470__A2 (.I(_08263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16471__B (.I(_07740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16478__A2 (.I(_08267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16487__A1 (.I(_08274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16491__A2 (.I(_08282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16491__B (.I(_08252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16495__B (.I(_08244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16497__A2 (.I(_08282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16497__B (.I(_08252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16503__B (.I(_08292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16504__A2 (.I(_08289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16508__B (.I(_08292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16509__A2 (.I(_08289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16514__B (.I(_08301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16515__A2 (.I(_08289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16520__A1 (.I(_08274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16521__A2 (.I(_08282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16521__B (.I(_08252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16525__A1 (.I(_08238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16526__A2 (.I(_08263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16527__I (.I(_01822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16528__B (.I(_08313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16530__A1 (.I(_08242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16531__A2 (.I(_08315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16533__A1 (.I(_08314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16534__I (.I(_07355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16535__A2 (.I(_08315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16535__B (.I(_08318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16536__A2 (.I(_08315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16542__A2 (.I(_08263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16543__B (.I(_08313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16548__A2 (.I(_08267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16551__A1 (.I(_08314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16557__A1 (.I(_08333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16558__I (.I(_01752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16559__A2 (.I(_08282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16559__B (.I(_08339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16563__B (.I(_08292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16566__B (.I(_08339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16571__B (.I(_08301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16573__A1 (.I(_08314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16576__B (.I(_08301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16578__A1 (.I(_08314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16582__B (.I(_08301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16584__A1 (.I(_08356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16588__A1 (.I(_08333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16589__B (.I(_08339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16593__A1 (.I(_08238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16594__A2 (.I(_08274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16595__B (.I(_08313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16596__A1 (.I(_08242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16599__A1 (.I(_08356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16600__A1 (.I(\tt_um_rejunity_sn76489.chan[1].attenuation.in ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16600__B (.I(_08318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16601__A1 (.I(\tt_um_rejunity_sn76489.chan[1].attenuation.in ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16602__A1 (.I(_01319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16603__I (.I(_08374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16605__A1 (.I(_01724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16605__A2 (.I(_08374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16609__A1 (.I(_01598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16611__A1 (.I(_01615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16612__I (.I(_08374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16613__I (.I(_08380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16615__I (.I(_08382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16618__A1 (.I(_01632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16620__I (.I(_08380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16621__I (.I(_08382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16624__A1 (.I(_01657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16626__I (.I(_08380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16627__I (.I(_08382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16628__A1 (.I(_01668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16631__A1 (.I(_01689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16632__I (.I(_08380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16633__I (.I(_08382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16636__A1 (.I(_01577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16637__A1 (.I(_01705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16638__A1 (.I(_01710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16639__A1 (.I(_01715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16646__A1 (.I(_08267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16647__A2 (.I(_08263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16648__B (.I(_08313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16653__A2 (.I(_08267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16656__A1 (.I(_08356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16661__A1 (.I(_08333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16662__B (.I(_08339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16666__B (.I(_08292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16668__B (.I(_01753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16674__A1 (.I(_08356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16675__I (.I(_06978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16679__A2 (.I(_08244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16680__A1 (.I(_08419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16684__A2 (.I(_08244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16685__A1 (.I(_08419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16689__A1 (.I(_08333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16690__A2 (.I(_08289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16690__B (.I(_01753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16694__A1 (.I(_08238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16695__A2 (.I(_08274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16696__B (.I(_01823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16697__A1 (.I(_08242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16698__A2 (.I(_08437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16700__A1 (.I(_08419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16701__A2 (.I(_08437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16701__B (.I(_08318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16702__A2 (.I(_08437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16706__A3 (.I(_03494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16708__I (.I(_08445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16709__I (.I(_08445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16710__B (.I(_08318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16711__A1 (.I(_03710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16712__I (.I(_01755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16716__A1 (.I(_08449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16718__I (.I(_08445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16720__A1 (.I(_08453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16723__A1 (.I(_08456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16725__A1 (.I(_01800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16727__B (.I(_08459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16728__A1 (.I(_01806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16732__I (.I(_08463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16733__I (.I(_08463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16734__B (.I(_08459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16735__A1 (.I(_03710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16736__B (.I(_08459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16737__A1 (.I(_08449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16738__I (.I(_08463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16739__B (.I(_08459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16740__A1 (.I(_08453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16743__A1 (.I(_08456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16745__A1 (.I(_01800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16747__A1 (.I(_01806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16749__I (.I(_00867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16750__I (.I(_00867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16752__A1 (.I(_03710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16755__A1 (.I(_08449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16756__I (.I(_00867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16758__A1 (.I(_08453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16760__A1 (.I(_08456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16762__A1 (.I(_01800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16763__I (.I(_02101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16764__B (.I(_00877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16765__A1 (.I(_01806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16766__I (.I(_03494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16768__A2 (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16772__I (.I(_00884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16773__I (.I(_00884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16774__A1 (.I(_03499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16775__C (.I(_02273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16776__A1 (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16777__I (.I(_02272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16779__A1 (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16781__A1 (.I(_02098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16787__I (.I(_00895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16788__I (.I(_00895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16789__A1 (.I(_03499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16792__A1 (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16794__C (.I(_00901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16795__A1 (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16796__C (.I(_00901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16797__A1 (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16798__C (.I(_00901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16799__A2 (.I(_01817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16801__I (.I(_00905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16802__I (.I(_00905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16803__A1 (.I(\tt_um_rejunity_sn76489.chan[1].attenuation.control[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16804__A1 (.I(_01741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16804__C (.I(_00901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16807__A1 (.I(_01756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16808__A1 (.I(\tt_um_rejunity_sn76489.chan[1].attenuation.control[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16809__A1 (.I(_08453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16811__A1 (.I(_08456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16812__B2 (.I(_01817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16814__I (.I(_00914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16815__I (.I(_00914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16817__A1 (.I(_01741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16820__A1 (.I(_01756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16822__A1 (.I(_01766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16824__A1 (.I(_01776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16827__A2 (.I(_04158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16828__A1 (.I(_00923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16828__B (.I(_01823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16831__C (.I(_07710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16833__C (.I(_04101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16834__C (.I(_04101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16836__A2 (.I(_03731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16836__B (.I(_00877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16838__A2 (.I(_03731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16839__A3 (.I(_03729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16840__A1 (.I(_06917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16842__B (.I(_01753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16844__B (.I(_00877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16848__A1 (.I(_08419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16849__A1 (.I(_01581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16849__A2 (.I(_03728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16850__I (.I(_00937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16851__I (.I(_00937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16852__C (.I(_01069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16853__A1 (.I(_02707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16854__A2 (.I(_02752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16855__A2 (.I(_03128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16855__A3 (.I(_03131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16857__A1 (.I(_02707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16857__A3 (.I(_03128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16857__A4 (.I(_02847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16865__A2 (.I(_02455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16865__B (.I(\channels.clk_div[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16866__A1 (.I(_03544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16866__A2 (.I(_03755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16866__A3 (.I(_00953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16869__A1 (.I(_00940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16874__B (.I(_00940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16878__A1 (.I(_00940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16881__I0 (.I(_00966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16881__S (.I(_00937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16891__A1 (.I(_01724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16891__A2 (.I(_00973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16893__S (.I(_00975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16895__S (.I(_00975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16897__I0 (.I(_00966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16897__S (.I(_00975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16899__S (.I(_00975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16913__A1 (.I(_03744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16913__A2 (.I(_03728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16913__B (.I(_01043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16915__S (.I(_00987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16917__S (.I(_00987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16919__I0 (.I(_00966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16919__S (.I(_00987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16921__S (.I(_00987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16926__A2 (.I(_00993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16926__B (.I(_00877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16927__A1 (.I(_01741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16927__A2 (.I(_00993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16928__A2 (.I(_00993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16928__B (.I(_02272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16929__A1 (.I(_08449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16929__A2 (.I(_00993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16930__A2 (.I(_00923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16931__A1 (.I(_01766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16931__A2 (.I(_00923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16958__CLK (.I(clknet_5_16__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16972__CLK (.I(clknet_5_23__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16991__CLK (.I(clknet_5_28__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__17016__CLK (.I(clknet_5_16__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__17030__CLK (.I(clknet_5_18__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__17048__CLK (.I(clknet_5_17__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__17055__D (.I(_00125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__17056__D (.I(_00126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__17057__D (.I(_00127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__17059__D (.I(_00129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__17128__CLK (.I(clknet_5_27__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__17162__CLK (.I(clknet_5_26__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__17208__CLK (.I(clknet_5_24__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__17237__CLK (.I(clknet_5_6__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__17240__CLK (.I(clknet_5_7__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__17250__CLK (.I(clknet_5_6__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__17319__D (.I(_00389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__17365__CLK (.I(clknet_5_25__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__17385__CLK (.I(clknet_5_31__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__17466__CLK (.I(clknet_5_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__17495__CLK (.I(clknet_5_5__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__17516__CLK (.I(clknet_5_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__17517__CLK (.I(clknet_5_2__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__17528__CLK (.I(clknet_5_6__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__17545__D (.I(_00615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__17547__D (.I(_00617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__17549__D (.I(_00619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__17563__CLK (.I(clknet_5_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__17564__CLK (.I(clknet_5_2__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__17572__CLK (.I(clknet_5_5__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__17572__D (.I(_00642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__17573__CLK (.I(clknet_5_5__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__17573__D (.I(_00643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__17574__D (.I(_00644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__17608__D (.I(_00678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__17635__CLK (.I(clknet_5_23__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__17638__CLK (.I(clknet_5_19__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__17667__D (.I(_00737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__17685__CLK (.I(clknet_5_11__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__17747__CLK (.I(clknet_5_8__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__17762__CLK (.I(clknet_5_9__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_0_clk_I (.I(clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_0_0_clk_I (.I(clknet_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_1_0_clk_I (.I(clknet_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_2_0_clk_I (.I(clknet_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_3_0_clk_I (.I(clknet_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_4_0_clk_I (.I(clknet_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_5_0_clk_I (.I(clknet_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_6_0_clk_I (.I(clknet_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_7_0_clk_I (.I(clknet_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_5_0__f_clk_I (.I(clknet_3_0_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_5_10__f_clk_I (.I(clknet_3_2_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_5_11__f_clk_I (.I(clknet_3_2_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_5_12__f_clk_I (.I(clknet_3_3_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_5_13__f_clk_I (.I(clknet_3_3_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_5_14__f_clk_I (.I(clknet_3_3_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_5_15__f_clk_I (.I(clknet_3_3_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_5_16__f_clk_I (.I(clknet_3_4_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_5_17__f_clk_I (.I(clknet_3_4_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_5_18__f_clk_I (.I(clknet_3_4_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_5_19__f_clk_I (.I(clknet_3_4_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_5_1__f_clk_I (.I(clknet_3_0_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_5_20__f_clk_I (.I(clknet_3_5_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_5_21__f_clk_I (.I(clknet_3_5_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_5_22__f_clk_I (.I(clknet_3_5_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_5_23__f_clk_I (.I(clknet_3_5_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_5_24__f_clk_I (.I(clknet_3_6_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_5_25__f_clk_I (.I(clknet_3_6_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_5_26__f_clk_I (.I(clknet_3_6_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_5_27__f_clk_I (.I(clknet_3_6_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_5_28__f_clk_I (.I(clknet_3_7_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_5_29__f_clk_I (.I(clknet_3_7_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_5_2__f_clk_I (.I(clknet_3_0_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_5_30__f_clk_I (.I(clknet_3_7_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_5_31__f_clk_I (.I(clknet_3_7_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_5_3__f_clk_I (.I(clknet_3_0_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_5_4__f_clk_I (.I(clknet_3_1_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_5_5__f_clk_I (.I(clknet_3_1_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_5_6__f_clk_I (.I(clknet_3_1_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_5_7__f_clk_I (.I(clknet_3_1_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_5_8__f_clk_I (.I(clknet_3_2_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_5_9__f_clk_I (.I(clknet_3_2_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_0_clk_I (.I(clknet_5_4__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_100_clk_I (.I(clknet_5_13__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_101_clk_I (.I(clknet_5_13__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_102_clk_I (.I(clknet_5_13__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_103_clk_I (.I(clknet_5_13__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_104_clk_I (.I(clknet_5_13__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_105_clk_I (.I(clknet_5_15__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_106_clk_I (.I(clknet_5_15__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_107_clk_I (.I(clknet_5_15__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_108_clk_I (.I(clknet_5_15__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_109_clk_I (.I(clknet_5_15__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_110_clk_I (.I(clknet_5_15__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_111_clk_I (.I(clknet_5_15__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_112_clk_I (.I(clknet_5_15__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_113_clk_I (.I(clknet_5_15__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_114_clk_I (.I(clknet_5_26__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_115_clk_I (.I(clknet_5_26__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_116_clk_I (.I(clknet_5_26__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_117_clk_I (.I(clknet_5_27__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_118_clk_I (.I(clknet_5_26__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_119_clk_I (.I(clknet_5_26__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_11_clk_I (.I(clknet_5_7__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_121_clk_I (.I(clknet_5_27__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_122_clk_I (.I(clknet_5_30__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_123_clk_I (.I(clknet_5_30__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_124_clk_I (.I(clknet_5_27__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_125_clk_I (.I(clknet_5_27__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_127_clk_I (.I(clknet_5_27__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_128_clk_I (.I(clknet_5_30__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_129_clk_I (.I(clknet_5_30__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_130_clk_I (.I(clknet_5_30__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_131_clk_I (.I(clknet_5_31__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_132_clk_I (.I(clknet_5_31__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_133_clk_I (.I(clknet_5_31__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_134_clk_I (.I(clknet_5_31__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_135_clk_I (.I(clknet_5_31__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_136_clk_I (.I(clknet_5_31__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_137_clk_I (.I(clknet_5_31__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_138_clk_I (.I(clknet_5_31__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_139_clk_I (.I(clknet_5_31__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_13_clk_I (.I(clknet_5_6__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_141_clk_I (.I(clknet_5_30__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_142_clk_I (.I(clknet_5_30__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_143_clk_I (.I(clknet_5_27__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_144_clk_I (.I(clknet_5_30__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_145_clk_I (.I(clknet_5_30__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_146_clk_I (.I(clknet_5_28__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_147_clk_I (.I(clknet_5_29__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_148_clk_I (.I(clknet_5_31__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_149_clk_I (.I(clknet_5_31__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_14_clk_I (.I(clknet_5_6__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_150_clk_I (.I(clknet_5_29__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_151_clk_I (.I(clknet_5_29__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_152_clk_I (.I(clknet_5_29__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_153_clk_I (.I(clknet_5_29__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_154_clk_I (.I(clknet_5_29__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_155_clk_I (.I(clknet_5_29__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_156_clk_I (.I(clknet_5_29__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_157_clk_I (.I(clknet_5_29__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_158_clk_I (.I(clknet_5_28__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_159_clk_I (.I(clknet_5_28__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_15_clk_I (.I(clknet_5_6__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_161_clk_I (.I(clknet_5_28__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_162_clk_I (.I(clknet_5_25__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_163_clk_I (.I(clknet_5_28__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_164_clk_I (.I(clknet_5_28__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_165_clk_I (.I(clknet_5_25__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_166_clk_I (.I(clknet_5_25__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_168_clk_I (.I(clknet_5_25__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_169_clk_I (.I(clknet_5_24__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_170_clk_I (.I(clknet_5_24__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_171_clk_I (.I(clknet_5_24__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_172_clk_I (.I(clknet_5_24__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_173_clk_I (.I(clknet_5_24__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_174_clk_I (.I(clknet_5_24__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_175_clk_I (.I(clknet_5_18__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_176_clk_I (.I(clknet_5_18__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_177_clk_I (.I(clknet_5_18__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_178_clk_I (.I(clknet_5_18__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_179_clk_I (.I(clknet_5_18__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_180_clk_I (.I(clknet_5_19__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_181_clk_I (.I(clknet_5_19__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_182_clk_I (.I(clknet_5_19__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_185_clk_I (.I(clknet_5_22__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_186_clk_I (.I(clknet_5_22__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_187_clk_I (.I(clknet_5_19__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_188_clk_I (.I(clknet_5_19__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_189_clk_I (.I(clknet_5_22__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_18_clk_I (.I(clknet_5_6__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_190_clk_I (.I(clknet_5_22__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_191_clk_I (.I(clknet_5_22__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_192_clk_I (.I(clknet_5_23__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_193_clk_I (.I(clknet_5_23__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_194_clk_I (.I(clknet_5_23__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_195_clk_I (.I(clknet_5_23__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_196_clk_I (.I(clknet_5_23__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_197_clk_I (.I(clknet_5_23__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_19_clk_I (.I(clknet_5_3__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_1_clk_I (.I(clknet_5_4__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_200_clk_I (.I(clknet_5_23__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_201_clk_I (.I(clknet_5_23__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_202_clk_I (.I(clknet_5_21__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_203_clk_I (.I(clknet_5_21__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_204_clk_I (.I(clknet_5_22__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_205_clk_I (.I(clknet_5_23__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_206_clk_I (.I(clknet_5_22__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_207_clk_I (.I(clknet_5_20__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_208_clk_I (.I(clknet_5_22__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_209_clk_I (.I(clknet_5_17__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_20_clk_I (.I(clknet_5_3__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_210_clk_I (.I(clknet_5_20__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_211_clk_I (.I(clknet_5_20__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_212_clk_I (.I(clknet_5_20__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_213_clk_I (.I(clknet_5_21__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_214_clk_I (.I(clknet_5_21__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_215_clk_I (.I(clknet_5_21__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_216_clk_I (.I(clknet_5_21__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_217_clk_I (.I(clknet_5_21__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_218_clk_I (.I(clknet_5_21__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_219_clk_I (.I(clknet_5_21__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_21_clk_I (.I(clknet_5_3__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_220_clk_I (.I(clknet_5_21__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_221_clk_I (.I(clknet_5_21__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_222_clk_I (.I(clknet_5_20__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_223_clk_I (.I(clknet_5_20__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_224_clk_I (.I(clknet_5_20__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_225_clk_I (.I(clknet_5_20__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_226_clk_I (.I(clknet_5_20__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_227_clk_I (.I(clknet_5_17__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_228_clk_I (.I(clknet_5_17__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_229_clk_I (.I(clknet_5_17__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_22_clk_I (.I(clknet_5_3__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_230_clk_I (.I(clknet_5_17__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_231_clk_I (.I(clknet_5_20__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_232_clk_I (.I(clknet_5_17__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_233_clk_I (.I(clknet_5_17__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_235_clk_I (.I(clknet_5_16__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_236_clk_I (.I(clknet_5_16__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_238_clk_I (.I(clknet_5_16__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_239_clk_I (.I(clknet_5_16__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_23_clk_I (.I(clknet_5_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_240_clk_I (.I(clknet_5_18__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_242_clk_I (.I(clknet_5_18__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_243_clk_I (.I(clknet_5_5__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_244_clk_I (.I(clknet_5_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_245_clk_I (.I(clknet_5_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_246_clk_I (.I(clknet_5_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_247_clk_I (.I(clknet_5_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_248_clk_I (.I(clknet_5_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_249_clk_I (.I(clknet_5_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_25_clk_I (.I(clknet_5_6__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_26_clk_I (.I(clknet_5_4__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_27_clk_I (.I(clknet_5_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_29_clk_I (.I(clknet_5_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_2_clk_I (.I(clknet_5_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_30_clk_I (.I(clknet_5_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_32_clk_I (.I(clknet_5_2__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_33_clk_I (.I(clknet_5_2__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_34_clk_I (.I(clknet_5_2__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_37_clk_I (.I(clknet_5_3__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_38_clk_I (.I(clknet_5_3__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_39_clk_I (.I(clknet_5_3__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_40_clk_I (.I(clknet_5_3__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_41_clk_I (.I(clknet_5_3__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_42_clk_I (.I(clknet_5_3__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_44_clk_I (.I(clknet_5_2__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_45_clk_I (.I(clknet_5_2__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_46_clk_I (.I(clknet_5_2__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_47_clk_I (.I(clknet_5_10__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_48_clk_I (.I(clknet_5_10__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_49_clk_I (.I(clknet_5_10__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_4_clk_I (.I(clknet_5_4__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_50_clk_I (.I(clknet_5_10__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_51_clk_I (.I(clknet_5_10__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_52_clk_I (.I(clknet_5_10__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_53_clk_I (.I(clknet_5_10__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_54_clk_I (.I(clknet_5_10__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_55_clk_I (.I(clknet_5_8__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_56_clk_I (.I(clknet_5_8__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_57_clk_I (.I(clknet_5_3__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_58_clk_I (.I(clknet_5_8__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_59_clk_I (.I(clknet_5_8__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_5_clk_I (.I(clknet_5_4__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_60_clk_I (.I(clknet_5_8__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_61_clk_I (.I(clknet_5_9__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_62_clk_I (.I(clknet_5_11__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_63_clk_I (.I(clknet_5_11__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_64_clk_I (.I(clknet_5_11__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_66_clk_I (.I(clknet_5_11__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_67_clk_I (.I(clknet_5_11__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_68_clk_I (.I(clknet_5_11__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_69_clk_I (.I(clknet_5_11__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_6_clk_I (.I(clknet_5_5__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_70_clk_I (.I(clknet_5_14__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_71_clk_I (.I(clknet_5_14__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_72_clk_I (.I(clknet_5_14__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_73_clk_I (.I(clknet_5_14__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_74_clk_I (.I(clknet_5_9__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_75_clk_I (.I(clknet_5_14__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_76_clk_I (.I(clknet_5_14__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_77_clk_I (.I(clknet_5_12__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_78_clk_I (.I(clknet_5_12__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_79_clk_I (.I(clknet_5_12__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_80_clk_I (.I(clknet_5_9__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_81_clk_I (.I(clknet_5_9__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_82_clk_I (.I(clknet_5_9__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_85_clk_I (.I(clknet_5_12__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_86_clk_I (.I(clknet_5_12__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_87_clk_I (.I(clknet_5_12__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_88_clk_I (.I(clknet_5_12__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_89_clk_I (.I(clknet_5_12__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_8_clk_I (.I(clknet_5_5__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_90_clk_I (.I(clknet_5_12__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_91_clk_I (.I(clknet_5_7__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_93_clk_I (.I(clknet_5_7__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_94_clk_I (.I(clknet_5_7__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_95_clk_I (.I(clknet_5_13__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_96_clk_I (.I(clknet_5_13__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_97_clk_I (.I(clknet_5_13__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_98_clk_I (.I(clknet_5_13__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_99_clk_I (.I(clknet_5_13__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_9_clk_I (.I(clknet_5_5__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input10_I (.I(bus_in[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input11_I (.I(bus_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input12_I (.I(bus_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input13_I (.I(bus_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input14_I (.I(bus_in[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input15_I (.I(bus_in[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input16_I (.I(bus_we));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input17_I (.I(rst));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1_I (.I(addr[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input2_I (.I(addr[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input3_I (.I(addr[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input4_I (.I(addr[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input5_I (.I(addr[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input6_I (.I(addr[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input7_I (.I(bus_cyc));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input8_I (.I(bus_in[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input9_I (.I(bus_in[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output19_I (.I(net19));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output20_I (.I(net20));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output22_I (.I(net22));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output23_I (.I(net23));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output25_I (.I(net25));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output26_I (.I(net26));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output27_I (.I(net27));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output28_I (.I(net28));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output29_I (.I(net29));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer10_I (.I(_05431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer11_I (.I(_05431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer19_I (.I(_05182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer20_I (.I(_05151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer28_I (.I(_04235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer31_I (.I(_04177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer6_I (.I(_05423_));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_100_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_100_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_100_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_100_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_100_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_100_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_100_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_100_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_100_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_100_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_100_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_100_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_100_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_100_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_100_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_100_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_101_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_101_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_101_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_101_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_101_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_101_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_101_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_101_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_101_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_101_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_101_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_101_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_102_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_102_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_102_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_102_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_102_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_102_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_102_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_102_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_102_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_102_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_102_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_102_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_102_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_102_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_102_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_102_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_103_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_103_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_103_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_103_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_103_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_103_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_103_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_103_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_103_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_103_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_103_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_103_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_103_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_104_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_104_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_104_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_104_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_104_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_104_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_104_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_104_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_104_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_104_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_104_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_105_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_105_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_105_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_105_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_105_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_105_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_105_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_105_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_105_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_105_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_105_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_105_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_106_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_106_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_106_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_106_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_106_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_106_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_106_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_106_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_106_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_106_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_106_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_106_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_106_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_106_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_107_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_107_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_107_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_107_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_107_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_107_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_107_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_107_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_107_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_107_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_107_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_107_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_108_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_108_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_108_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_108_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_108_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_109_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_109_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_109_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_109_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_109_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_109_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_109_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_10_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_10_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_10_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_10_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_110_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_110_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_110_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_110_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_110_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_110_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_110_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_110_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_110_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_110_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_110_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_111_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_111_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_111_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_111_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_111_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_111_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_111_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_112_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_112_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_112_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_112_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_112_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_112_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_112_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_112_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_112_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_112_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_112_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_113_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_113_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_113_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_113_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_113_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_113_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_113_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_113_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_113_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_113_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_113_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_113_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_113_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_114_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_114_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_114_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_114_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_114_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_114_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_114_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_114_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_114_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_114_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_114_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_114_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_114_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_114_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_114_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_114_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_115_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_115_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_115_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_115_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_115_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_115_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_115_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_115_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_115_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_115_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_116_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_116_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_116_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_116_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_116_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_116_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_116_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_116_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_116_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_116_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_116_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_116_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_116_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_116_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_116_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_116_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_116_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_117_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_117_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_117_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_117_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_117_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_117_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_117_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_117_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_117_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_117_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_117_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_117_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_117_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_118_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_118_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_118_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_118_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_118_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_118_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_118_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_118_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_118_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_118_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_118_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_118_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_118_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_118_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_119_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_119_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_119_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_119_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_119_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_119_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_119_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_119_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_119_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_11_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_11_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_11_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_11_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_11_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_11_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_11_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_120_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_120_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_120_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_120_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_120_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_120_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_120_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_120_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_120_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_120_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_120_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_120_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_121_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_121_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_121_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_121_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_121_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_121_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_121_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_121_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_121_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_122_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_122_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_122_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_122_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_122_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_122_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_122_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_122_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_122_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_122_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_122_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_122_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_122_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_122_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_123_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_123_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_123_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_123_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_123_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_123_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_123_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_123_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_123_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_123_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_123_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_123_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_123_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_124_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_124_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_124_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_124_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_124_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_124_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_124_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_124_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_124_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_124_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_124_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_124_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_124_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_124_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_124_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_125_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_125_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_125_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_125_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_125_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_125_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_125_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_125_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_125_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_125_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_125_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_125_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_126_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_126_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_126_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_126_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_126_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_126_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_126_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_126_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_126_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_126_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_126_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_126_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_126_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_126_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_127_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_127_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_127_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_127_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_127_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_127_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_127_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_127_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_127_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_127_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_127_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_127_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_127_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_127_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_128_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_128_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_128_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_128_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_128_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_128_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_128_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_128_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_128_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_128_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_128_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_128_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_128_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_128_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_129_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_129_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_129_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_129_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_129_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_129_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_129_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_129_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_129_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_129_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_129_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_129_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_129_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_129_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_129_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_129_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_129_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_129_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_129_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_129_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_129_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_129_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_129_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_129_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_12_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_12_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_12_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_12_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_130_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_130_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_130_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_130_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_130_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_130_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_130_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_130_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_130_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_130_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_130_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_130_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_130_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_130_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_130_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_130_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_130_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_130_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_130_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_130_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_130_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_131_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_131_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_131_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_131_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_131_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_131_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_131_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_132_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_132_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_132_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_132_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_132_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_133_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_133_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_133_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_133_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_133_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_133_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_133_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_133_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_133_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_133_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_133_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_133_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_133_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_133_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_133_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_133_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_133_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_133_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_133_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_133_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_133_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_133_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_134_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_134_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_134_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_134_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_134_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_134_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_134_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_134_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_134_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_135_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_135_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_135_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_135_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_135_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_135_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_135_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_135_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_135_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_135_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_136_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_136_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_136_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_136_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_136_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_136_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_136_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_136_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_136_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_136_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_136_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_136_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_136_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_136_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_136_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_136_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_136_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_137_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_137_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_137_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_137_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_137_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_137_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_137_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_137_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_137_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_137_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_137_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_137_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_138_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_138_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_138_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_138_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_138_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_138_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_138_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_138_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_138_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_139_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_139_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_139_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_139_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_139_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_139_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_139_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_139_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_139_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_139_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_139_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_139_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_139_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_139_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_139_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_139_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_139_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_139_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_139_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_139_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_139_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_139_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_139_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_13_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_13_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_13_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_13_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_13_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_13_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_13_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_13_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_140_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_140_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_140_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_140_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_140_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_140_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_140_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_140_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_140_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_140_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_140_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_140_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_140_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_140_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_140_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_140_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_140_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_140_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_140_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_140_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_140_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_140_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_140_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_141_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_141_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_141_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_141_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_141_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_141_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_141_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_141_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_141_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_141_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_141_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_141_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_141_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_141_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_141_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_141_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_141_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_141_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_141_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_141_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_141_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_141_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_141_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_141_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_141_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_141_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_142_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_142_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_142_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_142_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_142_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_142_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_142_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_142_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_142_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_142_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_142_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_142_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_142_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_142_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_142_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_142_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_142_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_142_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_142_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_142_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_142_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_142_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_142_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_143_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_143_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_143_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_143_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_143_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_143_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_143_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_143_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_143_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_143_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_143_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_143_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_143_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_143_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_143_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_143_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_143_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_143_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_143_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_143_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_143_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_143_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_143_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_143_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_143_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_144_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_144_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_144_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_144_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_144_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_144_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_144_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_144_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_144_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_144_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_144_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_144_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_144_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_144_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_144_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_144_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_144_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_144_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_145_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_145_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_145_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_145_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_145_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_145_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_145_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_145_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_145_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_145_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_145_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_145_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_145_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_145_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_145_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_145_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_145_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_145_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_145_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_145_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_145_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_145_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_145_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_145_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_146_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_146_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_146_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_146_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_146_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_146_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_146_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_146_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_146_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_146_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_146_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_146_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_146_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_146_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_146_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_146_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_146_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_146_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_146_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_146_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_146_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_146_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_146_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_146_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_146_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_146_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_146_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_147_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_147_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_147_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_147_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_147_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_147_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_147_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_147_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_147_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_147_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_147_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_147_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_147_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_147_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_147_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_147_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_147_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_147_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_147_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_147_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_147_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_147_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_147_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_147_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_147_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_147_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_147_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_147_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_147_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_147_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_147_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_148_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_148_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_148_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_148_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_148_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_148_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_148_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_148_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_148_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_148_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_148_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_148_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_148_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_148_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_148_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_148_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_148_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_148_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_148_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_148_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_148_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_148_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_148_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_148_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_148_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_148_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_148_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_148_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_148_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_149_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_149_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_149_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_149_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_149_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_149_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_149_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_149_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_149_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_149_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_149_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_149_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_149_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_149_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_149_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_149_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_149_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_149_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_149_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_149_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_149_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_149_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_149_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_149_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_149_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_149_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_149_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_149_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_149_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_149_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_14_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_14_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_14_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_14_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_14_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_14_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_14_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_150_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_150_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_150_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_150_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_150_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_150_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_150_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_150_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_150_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_150_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_150_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_150_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_150_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_150_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_150_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_150_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_150_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_150_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_150_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_150_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_150_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_150_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_150_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_150_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_151_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_151_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_151_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_151_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_151_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_151_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_151_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_151_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_151_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_151_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_151_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_151_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_151_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_151_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_151_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_151_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_151_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_151_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_151_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_151_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_151_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_151_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_151_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_152_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_152_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_152_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_152_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_152_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_152_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_152_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_152_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_152_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_152_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_152_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_152_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_152_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_152_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_152_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_152_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_152_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_152_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_152_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_152_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_152_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_152_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_153_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_153_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_153_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_153_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_153_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_153_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_153_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_153_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_153_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_153_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_153_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_153_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_153_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_153_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_153_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_153_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_153_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_153_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_154_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_154_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_154_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_154_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_154_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_154_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_154_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_154_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_154_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_154_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_154_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_154_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_154_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_154_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_154_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_154_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_154_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_154_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_154_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_154_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_154_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_154_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_154_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_155_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_155_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_155_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_155_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_155_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_155_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_155_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_155_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_155_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_155_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_155_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_155_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_155_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_155_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_155_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_155_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_155_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_155_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_155_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_155_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_155_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_155_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_155_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_155_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_155_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_156_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_156_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_156_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_156_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_156_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_156_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_156_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_156_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_156_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_156_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_156_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_156_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_156_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_156_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_156_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_156_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_156_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_156_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_156_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_156_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_156_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_156_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_156_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_156_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_156_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_156_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_156_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_156_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_156_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_156_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_156_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_156_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_156_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_156_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_156_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_156_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_156_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_156_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_156_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_156_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_156_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_156_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_156_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_156_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_156_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_156_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_156_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_156_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_156_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_156_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_156_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_156_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_157_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_157_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_157_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_157_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_157_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_157_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_157_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_157_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_157_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_157_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_157_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_157_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_157_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_157_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_157_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_157_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_157_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_157_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_157_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_157_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_157_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_157_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_157_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_157_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_157_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_157_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_157_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_157_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_157_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_157_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_157_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_157_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_157_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_157_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_157_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_157_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_157_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_157_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_157_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_157_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_157_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_157_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_157_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_157_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_157_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_157_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_157_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_157_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_157_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_157_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_157_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_157_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_157_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_157_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_157_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_157_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_158_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_158_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_158_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_158_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_158_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_158_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_158_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_158_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_158_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_158_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_158_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_158_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_158_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_158_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_158_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_158_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_158_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_158_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_158_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_158_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_158_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_158_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_158_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_158_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_158_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_158_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_158_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_158_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_158_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_158_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_158_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_158_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_158_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_158_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_158_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_158_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_158_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_158_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_158_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_158_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_158_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_158_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_158_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_158_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_158_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_158_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_158_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_158_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_158_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_158_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_158_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_159_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_159_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_159_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_159_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_159_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_159_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_159_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_159_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_159_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_159_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_159_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_159_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_159_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_159_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_159_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_159_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_159_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_159_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_159_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_159_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_159_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_159_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_159_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_159_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_159_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_159_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_159_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_159_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_159_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_159_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_159_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_159_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_159_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_159_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_159_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_159_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_159_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_159_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_159_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_159_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_159_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_159_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_159_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_159_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_159_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_159_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_159_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_15_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_160_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_160_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_160_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_160_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_160_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_160_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_160_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_160_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_160_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_160_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_160_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_160_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_160_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_160_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_160_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_160_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_160_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_160_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_160_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_160_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_160_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_160_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_160_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_160_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_160_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_160_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_160_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_160_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_160_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_160_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_160_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_160_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_160_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_160_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_160_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_160_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_160_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_160_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_160_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_160_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_160_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_160_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_160_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_160_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_160_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_160_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_160_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_160_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_160_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_160_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_160_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_160_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_160_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_160_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_160_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_160_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_160_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_160_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_160_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_160_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_161_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_161_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_161_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_161_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_161_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_161_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_161_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_161_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_161_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_161_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_161_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_161_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_161_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_161_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_161_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_161_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_161_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_161_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_161_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_161_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_161_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_161_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_161_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_161_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_161_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_161_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_161_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_161_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_161_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_161_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_161_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_161_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_161_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_161_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_161_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_161_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_161_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_161_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_161_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_161_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_161_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_161_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_161_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_161_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_161_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_162_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_162_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_162_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_162_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_162_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_162_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_162_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_162_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_162_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_162_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_162_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_162_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_162_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_162_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_162_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_162_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_162_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_162_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_162_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_162_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_162_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_162_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_162_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_162_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_162_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_162_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_162_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_162_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_162_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_162_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_162_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_162_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_162_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_162_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_162_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_162_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_162_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_162_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_162_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_162_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_162_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_162_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_162_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_162_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_162_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_162_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_162_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_162_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_162_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_163_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_163_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_163_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_163_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_163_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_163_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_163_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_163_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_163_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_163_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_163_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_163_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_163_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_163_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_163_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_163_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_163_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_163_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_163_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_163_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_163_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_163_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_163_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_163_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_163_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_163_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_163_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_163_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_163_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_163_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_163_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_163_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_163_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_163_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_163_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_163_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_163_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_163_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_163_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_163_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_163_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_163_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_163_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_163_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_163_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_163_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_163_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_163_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_163_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_163_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_163_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_163_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_163_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_163_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_164_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_164_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_164_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_164_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_164_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_164_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_164_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_164_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_164_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_164_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_164_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_164_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_164_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_164_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_164_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_164_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_164_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_164_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_164_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_164_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_164_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_164_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_164_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_164_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_164_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_164_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_164_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_164_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_164_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_164_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_164_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_164_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_164_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_164_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_164_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_164_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_164_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_164_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_164_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_164_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_164_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_164_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_164_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_164_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_164_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_164_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_164_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_164_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_164_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_164_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_164_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_164_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_164_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_164_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_164_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_164_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_164_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_164_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_164_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_164_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_164_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_164_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_165_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_165_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_165_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_165_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_165_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_165_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_165_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_165_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_165_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_165_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_165_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_165_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_165_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_165_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_165_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_165_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_165_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_165_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_165_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_165_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_165_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_165_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_165_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_165_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_165_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_165_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_165_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_165_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_165_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_165_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_165_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_165_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_165_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_165_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_165_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_165_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_165_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_165_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_165_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_165_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_165_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_165_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_165_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_165_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_165_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_165_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_165_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_165_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_165_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_165_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_165_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_165_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_165_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_165_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_165_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_165_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_165_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_165_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_165_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_165_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_165_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_165_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_165_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_165_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_165_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_165_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_165_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_165_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_165_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_165_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_165_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_165_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_165_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_165_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_165_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_165_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_165_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_165_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_165_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_165_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_166_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_166_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_166_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_166_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_166_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_166_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_166_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_166_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_166_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_166_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_166_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_166_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_166_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_166_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_166_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_166_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_166_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_166_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_166_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_166_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_166_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_166_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_166_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_166_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_166_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_166_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_166_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_166_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_166_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_166_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_166_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_166_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_166_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_166_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_166_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_166_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_166_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_166_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_166_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_166_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_166_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_166_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_166_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_166_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_166_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_166_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_166_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_166_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_166_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_166_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_166_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_166_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_166_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_166_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_166_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_166_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_166_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_166_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_166_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_166_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_166_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_166_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_166_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_166_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_166_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_166_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_166_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_166_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_166_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_166_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_166_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_166_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_166_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_166_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_166_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_166_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_166_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_166_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_166_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_166_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_166_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_166_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_166_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_166_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_167_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_167_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_167_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_167_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_167_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_167_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_167_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_167_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_167_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_167_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_167_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_167_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_167_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_167_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_167_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_167_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_167_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_167_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_167_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_167_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_167_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_167_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_167_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_167_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_167_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_167_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_167_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_167_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_167_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_167_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_167_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_167_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_167_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_167_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_167_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_167_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_167_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_167_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_167_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_167_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_167_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_167_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_167_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_167_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_167_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_167_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_167_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_167_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_167_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_167_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_167_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_167_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_167_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_167_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_167_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_167_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_167_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_167_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_167_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_167_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_167_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_167_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_167_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_167_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_167_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_167_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_167_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_167_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_167_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_167_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_167_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_167_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_167_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_167_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_167_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_167_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_167_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_167_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_167_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_167_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_167_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_167_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_167_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_167_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_167_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_167_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_167_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_167_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_167_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_167_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_167_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_167_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_167_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_168_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_168_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_168_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_168_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_168_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_168_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_168_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_168_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_168_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_168_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_168_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_168_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_168_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_168_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_168_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_168_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_168_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_168_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_168_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_168_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_168_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_168_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_168_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_168_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_168_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_168_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_168_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_168_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_168_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_168_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_168_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_168_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_168_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_168_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_168_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_168_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_168_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_168_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_168_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_168_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_168_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_168_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_168_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_168_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_168_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_168_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_168_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_168_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_168_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_168_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_168_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_168_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_168_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_168_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_168_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_168_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_168_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_168_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_168_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_168_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_168_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_168_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_168_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_168_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_168_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_168_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_168_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_168_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_168_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_168_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_168_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_168_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_168_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_168_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_168_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_168_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_168_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_168_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_168_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_168_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_168_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_168_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_168_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_168_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_168_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_168_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_168_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_169_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_169_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_169_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_169_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_169_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_169_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_169_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_169_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_169_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_169_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_169_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_169_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_169_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_169_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_169_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_169_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_169_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_16_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_16_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_16_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_16_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_16_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_170_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_170_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_170_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_170_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_170_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_170_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_170_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_170_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_170_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_170_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_170_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_170_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_170_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_170_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_170_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_170_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_170_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_170_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_170_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_170_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_170_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_170_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_170_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_170_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_170_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_170_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_170_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_170_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_170_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_170_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_170_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_170_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_170_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_170_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_170_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_170_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_170_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_170_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_170_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_170_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_170_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_170_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_170_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_170_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_170_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_170_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_170_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_170_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_170_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_170_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_170_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_170_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_170_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_170_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_170_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_170_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_170_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_170_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_170_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_170_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_170_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_170_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_170_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_170_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_170_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_170_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_170_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_170_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_170_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_170_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_170_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_170_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_170_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_170_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_170_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_170_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_170_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_170_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_170_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_170_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_170_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_170_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_170_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_170_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_170_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_170_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_170_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_170_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_170_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_170_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_170_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_170_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_170_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_170_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_170_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_170_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_170_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_170_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_170_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_170_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_170_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_170_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_170_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_170_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_170_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_170_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_170_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_171_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_171_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_171_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_171_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_171_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_171_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_171_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_171_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_171_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_171_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_171_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_171_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_171_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_171_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_171_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_171_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_171_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_171_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_171_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_171_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_171_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_171_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_171_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_171_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_171_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_171_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_171_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_171_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_171_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_171_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_171_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_171_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_171_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_171_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_171_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_171_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_171_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_171_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_171_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_171_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_171_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_171_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_171_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_171_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_171_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_171_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_171_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_171_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_171_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_171_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_171_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_171_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_171_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_171_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_171_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_171_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_171_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_171_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_171_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_171_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_171_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_171_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_171_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_171_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_171_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_171_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_171_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_171_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_171_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_171_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_171_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_171_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_171_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_171_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_171_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_172_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_172_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_172_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_172_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_172_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_172_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_172_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_172_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_172_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_172_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_172_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_172_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_172_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_172_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_172_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_172_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_172_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_172_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_172_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_172_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_172_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_172_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_172_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_172_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_172_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_172_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_172_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_172_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_172_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_172_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_172_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_172_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_172_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_172_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_172_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_172_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_172_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_172_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_172_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_172_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_172_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_172_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_172_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_172_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_172_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_172_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_172_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_172_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_172_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_172_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_172_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_172_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_172_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_172_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_172_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_172_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_172_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_172_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_172_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_172_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_172_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_172_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_172_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_172_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_172_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_172_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_172_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_172_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_172_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_172_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_172_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_172_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_172_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_172_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_172_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_172_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_172_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_172_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_172_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_172_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_172_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_172_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_172_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_172_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_172_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_172_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_172_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_172_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_173_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_173_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_173_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_173_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_173_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_173_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_173_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_173_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_173_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_173_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_173_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_173_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_173_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_173_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_173_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_173_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_173_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_173_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_173_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_173_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_173_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_173_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_173_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_173_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_173_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_173_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_173_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_173_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_173_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_173_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_173_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_173_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_173_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_173_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_173_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_173_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_173_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_173_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_173_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_173_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_173_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_173_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_173_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_173_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_173_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_173_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_173_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_173_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_173_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_173_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_173_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_173_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_173_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_173_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_173_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_173_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_173_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_173_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_173_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_173_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_173_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_173_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_173_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_173_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_173_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_173_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_173_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_173_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_173_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_173_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_173_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_173_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_173_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_173_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_173_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_173_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_173_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_173_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_173_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_173_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_173_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_173_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_173_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_174_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_174_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_174_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_174_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_174_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_174_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_174_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_174_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_174_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_174_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_174_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_174_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_174_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_174_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_174_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_174_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_174_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_174_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_174_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_174_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_174_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_174_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_174_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_174_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_174_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_174_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_174_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_174_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_174_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_174_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_174_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_174_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_174_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_174_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_174_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_174_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_174_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_174_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_174_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_174_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_174_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_174_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_174_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_174_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_174_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_174_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_174_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_174_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_174_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_174_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_174_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_174_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_174_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_174_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_174_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_174_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_174_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_174_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_174_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_174_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_174_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_174_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_174_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_174_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_174_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_174_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_174_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_174_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_174_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_174_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_174_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_174_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_174_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_174_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_174_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_174_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_174_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_174_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_174_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_174_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_174_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_174_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_174_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_174_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_174_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_174_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_174_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_174_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_174_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_174_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_174_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_174_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_174_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_174_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_174_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_174_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_174_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_174_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_174_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_174_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_174_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_174_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_174_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_174_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_174_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_174_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_174_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_174_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_174_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_174_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_174_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_174_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_174_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_174_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_174_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_174_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_174_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_174_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_174_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_174_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_175_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_175_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_175_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_175_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_175_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_175_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_175_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_175_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_175_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_175_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_175_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_175_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_175_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_175_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_175_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_175_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_175_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_175_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_175_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_175_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_175_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_175_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_175_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_175_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_175_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_175_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_175_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_175_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_175_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_175_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_175_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_175_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_175_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_175_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_175_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_175_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_175_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_175_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_175_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_175_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_175_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_175_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_175_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_175_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_175_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_175_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_175_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_175_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_175_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_175_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_175_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_175_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_175_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_175_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_175_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_175_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_175_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_175_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_175_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_175_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_175_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_175_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_175_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_175_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_175_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_175_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_175_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_175_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_175_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_175_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_175_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_175_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_175_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_175_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_175_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_175_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_175_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_175_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_175_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_175_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_175_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_175_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_175_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_175_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_175_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_175_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_175_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_175_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_175_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_175_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_175_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_175_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_175_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_175_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_175_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_175_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_175_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_176_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_176_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_176_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_176_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_176_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_176_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_176_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_176_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_176_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_176_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_176_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_176_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_176_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_176_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_176_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_176_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_176_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_176_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_176_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_176_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_176_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_176_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_176_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_176_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_176_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_176_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_176_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_176_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_176_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_176_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_176_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_176_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_176_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_176_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_176_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_176_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_176_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_176_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_176_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_176_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_176_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_176_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_176_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_176_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_176_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_176_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_176_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_176_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_176_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_176_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_176_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_176_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_176_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_176_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_176_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_176_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_176_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_176_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_176_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_176_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_176_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_176_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_176_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_176_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_176_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_176_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_176_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_176_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_176_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_176_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_176_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_176_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_176_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_176_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_176_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_176_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_176_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_176_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_176_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_176_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_176_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_176_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_176_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_176_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_176_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_176_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_176_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_176_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_176_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_176_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_176_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_176_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_176_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_176_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_176_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_176_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_176_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_176_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_176_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_176_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_176_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_176_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_176_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_176_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_176_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_176_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_176_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_176_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_176_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_176_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_176_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_176_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_176_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_176_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_177_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_177_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_177_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_177_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_177_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_177_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_177_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_177_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_177_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_177_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_177_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_177_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_177_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_177_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_177_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_177_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_177_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_177_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_177_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_177_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_177_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_177_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_177_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_177_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_177_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_177_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_177_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_177_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_177_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_177_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_177_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_177_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_177_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_177_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_177_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_177_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_177_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_177_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_177_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_177_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_177_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_177_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_177_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_177_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_177_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_177_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_177_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_177_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_177_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_177_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_177_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_177_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_177_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_177_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_177_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_177_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_177_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_177_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_177_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_177_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_177_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_177_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_177_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_177_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_177_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_177_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_177_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_177_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_177_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_177_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_177_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_177_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_177_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_177_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_177_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_177_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_177_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_177_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_177_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_177_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_177_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_177_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_177_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_177_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_177_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_177_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_177_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_177_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_177_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_177_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_177_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_177_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_177_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_177_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_177_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_177_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_177_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_177_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_177_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_177_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_178_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_178_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_178_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_178_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_178_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_178_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_178_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_178_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_178_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_178_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_178_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_178_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_178_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_178_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_178_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_178_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_178_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_178_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_178_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_178_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_178_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_178_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_178_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_178_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_178_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_178_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_178_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_178_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_178_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_178_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_178_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_178_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_178_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_178_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_178_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_178_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_178_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_178_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_178_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_178_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_178_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_178_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_178_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_178_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_178_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_178_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_178_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_178_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_178_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_178_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_178_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_178_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_178_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_178_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_178_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_178_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_178_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_178_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_178_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_178_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_178_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_178_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_178_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_178_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_178_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_178_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_178_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_178_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_178_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_178_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_178_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_178_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_178_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_178_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_178_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_178_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_178_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_178_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_178_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_178_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_178_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_178_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_178_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_178_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_178_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_178_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_178_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_178_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_178_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_178_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_178_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_178_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_178_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_178_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_178_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_178_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_178_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_178_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_178_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_178_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_178_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_178_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_178_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_178_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_178_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_178_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_178_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_178_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_178_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_178_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_179_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_179_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_179_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_179_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_179_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_179_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_179_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_179_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_179_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_179_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_179_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_179_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_179_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_179_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_179_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_179_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_179_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_179_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_179_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_179_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_179_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_179_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_179_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_179_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_179_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_179_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_179_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_179_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_179_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_179_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_179_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_179_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_179_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_179_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_179_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_179_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_179_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_179_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_179_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_179_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_179_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_179_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_179_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_179_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_179_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_179_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_179_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_179_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_179_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_179_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_179_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_179_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_179_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_179_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_179_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_179_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_179_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_179_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_179_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_179_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_179_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_179_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_179_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_179_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_179_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_179_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_179_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_179_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_179_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_179_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_179_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_179_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_179_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_179_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_179_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_179_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_179_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_179_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_179_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_179_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_179_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_179_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_179_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_179_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_179_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_179_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_179_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_179_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_179_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_179_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_179_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_179_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_179_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_17_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_17_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_17_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_180_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_180_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_180_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_180_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_180_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_180_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_180_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_180_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_180_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_180_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_180_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_180_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_180_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_180_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_180_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_180_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_180_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_180_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_180_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_180_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_180_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_180_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_180_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_180_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_180_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_180_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_180_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_180_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_180_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_180_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_180_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_180_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_180_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_180_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_180_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_180_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_180_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_180_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_180_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_180_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_180_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_180_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_180_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_180_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_180_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_180_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_180_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_180_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_180_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_180_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_180_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_180_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_180_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_180_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_180_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_180_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_180_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_180_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_180_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_180_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_180_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_180_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_180_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_180_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_180_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_180_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_180_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_180_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_180_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_180_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_180_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_180_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_180_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_180_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_180_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_180_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_180_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_180_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_180_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_181_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_181_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_181_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_181_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_181_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_181_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_181_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_181_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_181_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_181_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_181_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_181_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_181_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_181_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_181_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_181_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_181_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_181_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_181_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_181_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_181_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_181_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_181_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_181_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_181_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_181_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_181_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_181_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_181_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_181_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_181_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_181_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_181_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_181_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_181_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_181_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_181_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_181_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_181_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_181_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_181_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_181_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_181_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_181_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_181_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_181_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_181_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_181_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_181_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_181_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_181_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_181_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_181_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_181_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_181_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_181_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_181_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_181_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_181_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_181_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_181_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_181_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_181_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_181_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_181_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_181_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_181_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_181_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_181_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_181_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_181_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_181_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_181_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_181_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_181_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_181_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_181_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_181_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_181_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_181_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_181_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_181_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_181_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_181_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_181_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_181_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_181_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_181_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_181_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_182_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_182_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_182_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_182_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_182_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_182_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_182_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_182_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_182_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_182_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_182_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_182_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_182_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_182_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_182_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_182_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_182_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_182_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_182_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_182_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_182_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_182_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_182_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_182_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_182_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_182_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_182_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_182_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_182_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_182_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_182_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_182_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_182_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_182_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_182_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_182_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_182_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_182_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_182_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_182_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_182_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_182_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_182_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_182_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_182_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_182_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_182_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_182_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_182_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_182_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_182_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_182_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_182_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_182_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_182_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_182_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_182_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_182_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_182_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_182_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_182_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_182_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_182_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_182_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_182_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_182_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_182_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_182_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_182_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_182_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_182_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_182_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_182_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_182_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_182_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_182_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_182_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_182_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_182_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_182_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_182_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_182_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_182_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_182_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_182_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_182_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_182_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_182_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_182_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_182_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_182_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_182_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_182_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_182_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_182_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_182_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_182_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_182_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_182_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_182_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_182_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_182_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_182_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_182_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_182_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_182_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_182_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_182_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_182_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_182_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_182_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_18_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_18_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_18_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_19_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_19_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_19_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_20_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_20_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_20_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_21_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_21_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_22_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_22_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_22_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_22_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_22_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_23_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_23_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_23_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_24_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_24_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_24_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_25_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_25_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_25_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_25_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_26_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_26_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_26_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_27_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_27_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_27_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_27_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_28_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_28_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_29_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_29_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_29_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_29_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_29_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_30_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_30_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_31_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_32_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_32_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_33_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_33_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_33_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_33_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_34_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_34_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_34_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_35_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_35_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_35_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_36_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_36_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_37_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_39_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_39_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_39_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_39_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_39_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_39_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_3_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_3_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_3_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_3_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_3_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_3_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_3_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_3_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_3_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_40_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_40_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_40_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_40_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_40_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_40_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_41_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_41_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_41_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_41_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_42_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_42_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_43_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_43_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_44_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_44_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_45_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_45_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_45_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_45_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_46_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_46_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_46_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_46_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_46_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_48_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_48_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_49_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_49_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_49_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_49_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_4_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_4_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_50_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_50_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_50_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_50_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_50_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_51_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_51_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_51_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_51_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_51_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_51_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_52_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_52_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_53_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_53_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_53_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_53_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_54_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_54_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_54_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_55_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_55_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_56_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_56_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_56_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_57_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_57_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_57_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_58_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_58_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_58_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_59_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_59_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_59_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_59_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_5_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_5_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_5_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_5_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_5_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_5_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_60_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_60_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_60_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_61_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_61_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_61_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_62_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_63_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_63_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_64_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_64_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_64_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_65_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_65_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_66_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_67_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_67_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_67_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_67_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_67_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_68_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_68_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_68_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_68_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_68_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_68_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_68_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_69_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_69_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_6_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_6_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_6_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_6_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_6_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_6_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_6_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_6_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_70_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_71_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_71_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_71_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_72_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_72_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_72_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_72_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_73_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_73_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_73_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_73_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_74_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_74_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_75_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_76_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_76_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_76_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_76_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_77_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_77_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_77_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_78_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_78_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_78_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_78_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_78_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_78_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_78_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_79_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_79_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_79_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_79_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_7_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_7_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_7_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_7_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_7_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_80_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_80_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_81_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_81_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_82_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_82_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_83_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_83_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_83_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_83_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_83_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_83_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_83_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_83_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_83_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_83_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_83_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_84_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_84_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_84_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_84_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_84_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_84_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_84_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_84_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_84_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_84_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_84_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_84_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_84_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_85_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_85_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_85_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_85_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_85_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_85_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_85_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_85_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_85_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_85_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_85_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_85_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_85_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_85_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_86_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_86_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_86_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_86_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_86_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_86_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_86_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_86_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_86_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_87_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_87_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_87_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_87_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_87_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_87_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_87_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_88_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_89_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_89_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_89_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_89_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_8_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_8_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_8_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_90_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_90_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_90_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_90_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_90_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_90_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_91_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_91_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_91_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_91_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_91_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_91_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_91_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_91_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_91_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_91_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_91_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_92_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_93_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_93_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_93_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_93_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_93_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_93_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_93_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_93_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_93_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_93_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_93_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_94_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_94_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_94_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_94_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_94_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_94_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_94_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_94_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_94_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_94_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_94_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_95_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_95_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_95_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_95_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_95_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_95_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_95_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_95_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_95_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_95_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_95_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_95_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_95_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_96_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_96_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_96_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_96_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_96_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_96_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_96_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_96_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_96_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_97_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_97_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_97_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_97_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_97_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_97_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_97_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_97_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_97_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_97_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_97_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_98_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_98_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_98_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_98_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_98_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_98_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_98_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_98_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_98_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_98_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_98_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_98_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_98_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_99_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_99_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_99_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_99_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_99_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_99_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_99_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_9_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_9_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_9_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_979 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_Left_183 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_Right_0 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_100_Left_283 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_100_Right_100 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_101_Left_284 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_101_Right_101 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_102_Left_285 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_102_Right_102 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_103_Left_286 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_103_Right_103 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_104_Left_287 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_104_Right_104 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_105_Left_288 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_105_Right_105 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_106_Left_289 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_106_Right_106 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_107_Left_290 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_107_Right_107 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_108_Left_291 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_108_Right_108 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_109_Left_292 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_109_Right_109 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_Left_193 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_Right_10 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_110_Left_293 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_110_Right_110 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_111_Left_294 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_111_Right_111 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_112_Left_295 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_112_Right_112 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_113_Left_296 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_113_Right_113 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_114_Left_297 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_114_Right_114 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_115_Left_298 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_115_Right_115 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_116_Left_299 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_116_Right_116 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_117_Left_300 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_117_Right_117 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_118_Left_301 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_118_Right_118 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_119_Left_302 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_119_Right_119 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_Left_194 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_Right_11 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_120_Left_303 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_120_Right_120 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_121_Left_304 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_121_Right_121 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_122_Left_305 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_122_Right_122 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_123_Left_306 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_123_Right_123 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_124_Left_307 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_124_Right_124 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_125_Left_308 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_125_Right_125 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_126_Left_309 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_126_Right_126 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_127_Left_310 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_127_Right_127 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_128_Left_311 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_128_Right_128 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_129_Left_312 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_129_Right_129 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_Left_195 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_Right_12 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_130_Left_313 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_130_Right_130 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_131_Left_314 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_131_Right_131 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_132_Left_315 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_132_Right_132 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_133_Left_316 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_133_Right_133 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_134_Left_317 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_134_Right_134 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_135_Left_318 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_135_Right_135 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_136_Left_319 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_136_Right_136 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_137_Left_320 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_137_Right_137 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_138_Left_321 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_138_Right_138 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_139_Left_322 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_139_Right_139 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_Left_196 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_Right_13 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_140_Left_323 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_140_Right_140 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_141_Left_324 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_141_Right_141 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_142_Left_325 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_142_Right_142 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_143_Left_326 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_143_Right_143 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_144_Left_327 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_144_Right_144 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_145_Left_328 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_145_Right_145 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_146_Left_329 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_146_Right_146 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_147_Left_330 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_147_Right_147 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_148_Left_331 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_148_Right_148 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_149_Left_332 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_149_Right_149 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_Left_197 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_Right_14 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_150_Left_333 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_150_Right_150 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_151_Left_334 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_151_Right_151 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_152_Left_335 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_152_Right_152 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_153_Left_336 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_153_Right_153 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_154_Left_337 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_154_Right_154 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_155_Left_338 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_155_Right_155 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_156_Left_339 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_156_Right_156 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_157_Left_340 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_157_Right_157 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_158_Left_341 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_158_Right_158 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_159_Left_342 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_159_Right_159 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_Left_198 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_Right_15 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_160_Left_343 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_160_Right_160 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_161_Left_344 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_161_Right_161 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_162_Left_345 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_162_Right_162 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_163_Left_346 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_163_Right_163 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_164_Left_347 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_164_Right_164 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_165_Left_348 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_165_Right_165 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_166_Left_349 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_166_Right_166 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_167_Left_350 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_167_Right_167 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_168_Left_351 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_168_Right_168 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_169_Left_352 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_169_Right_169 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_Left_199 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_Right_16 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_170_Left_353 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_170_Right_170 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_171_Left_354 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_171_Right_171 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_172_Left_355 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_172_Right_172 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_173_Left_356 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_173_Right_173 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_174_Left_357 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_174_Right_174 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_175_Left_358 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_175_Right_175 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_176_Left_359 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_176_Right_176 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_177_Left_360 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_177_Right_177 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_178_Left_361 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_178_Right_178 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_179_Left_362 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_179_Right_179 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_Left_200 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_Right_17 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_180_Left_363 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_180_Right_180 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_181_Left_364 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_181_Right_181 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_182_Left_365 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_182_Right_182 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_Left_201 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_Right_18 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_Left_202 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_Right_19 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_Left_184 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_Right_1 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_Left_203 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_Right_20 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_Left_204 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_Right_21 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_Left_205 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_Right_22 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_Left_206 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_Right_23 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_Left_207 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_Right_24 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_Left_208 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_Right_25 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_Left_209 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_Right_26 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_Left_210 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_Right_27 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_Left_211 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_Right_28 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_Left_212 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_Right_29 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_Left_185 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_Right_2 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_Left_213 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_Right_30 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_Left_214 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_Right_31 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_Left_215 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_Right_32 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_Left_216 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_Right_33 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_Left_217 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_Right_34 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_Left_218 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_Right_35 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_Left_219 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_Right_36 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_Left_220 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_Right_37 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_Left_221 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_Right_38 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_Left_222 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_Right_39 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_Left_186 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_Right_3 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_Left_223 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_Right_40 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_Left_224 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_Right_41 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_Left_225 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_Right_42 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_Left_226 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_Right_43 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_Left_227 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_Right_44 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_Left_228 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_Right_45 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_Left_229 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_Right_46 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_47_Left_230 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_47_Right_47 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_48_Left_231 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_48_Right_48 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_49_Left_232 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_49_Right_49 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_Left_187 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_Right_4 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_50_Left_233 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_50_Right_50 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_51_Left_234 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_51_Right_51 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_52_Left_235 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_52_Right_52 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_53_Left_236 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_53_Right_53 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_54_Left_237 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_54_Right_54 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_55_Left_238 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_55_Right_55 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_56_Left_239 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_56_Right_56 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_57_Left_240 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_57_Right_57 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_58_Left_241 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_58_Right_58 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_59_Left_242 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_59_Right_59 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_Left_188 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_Right_5 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_60_Left_243 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_60_Right_60 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_61_Left_244 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_61_Right_61 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_62_Left_245 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_62_Right_62 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_63_Left_246 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_63_Right_63 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_64_Left_247 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_64_Right_64 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_65_Left_248 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_65_Right_65 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_66_Left_249 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_66_Right_66 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_67_Left_250 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_67_Right_67 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_68_Left_251 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_68_Right_68 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_69_Left_252 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_69_Right_69 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_Left_189 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_Right_6 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_70_Left_253 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_70_Right_70 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_71_Left_254 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_71_Right_71 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_72_Left_255 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_72_Right_72 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_73_Left_256 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_73_Right_73 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_74_Left_257 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_74_Right_74 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_75_Left_258 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_75_Right_75 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_76_Left_259 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_76_Right_76 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_77_Left_260 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_77_Right_77 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_78_Left_261 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_78_Right_78 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_79_Left_262 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_79_Right_79 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_Left_190 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_Right_7 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_80_Left_263 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_80_Right_80 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_81_Left_264 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_81_Right_81 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_82_Left_265 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_82_Right_82 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_83_Left_266 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_83_Right_83 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_84_Left_267 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_84_Right_84 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_85_Left_268 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_85_Right_85 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_86_Left_269 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_86_Right_86 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_87_Left_270 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_87_Right_87 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_88_Left_271 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_88_Right_88 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_89_Left_272 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_89_Right_89 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_Left_191 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_Right_8 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_90_Left_273 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_90_Right_90 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_91_Left_274 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_91_Right_91 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_92_Left_275 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_92_Right_92 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_93_Left_276 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_93_Right_93 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_94_Left_277 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_94_Right_94 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_95_Left_278 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_95_Right_95 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_96_Left_279 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_96_Right_96 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_97_Left_280 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_97_Right_97 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_98_Left_281 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_98_Right_98 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_99_Left_282 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_99_Right_99 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_Left_192 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_Right_9 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_2254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_2255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_2256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_2257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_2258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_2259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_2260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_2261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_2262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_2263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_2264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_2265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_2266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_2268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_2269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_2270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_2272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_2275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_2276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_2277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_2278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_2279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_2280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_2281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_2282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_2283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_2284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_2285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_2286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_2287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_2288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_2289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_2290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_2291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_2292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_2293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_2294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_2295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_2296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_2297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_2298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_2299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_2300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_2301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_2303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_2304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_2305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_2307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_2308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_2310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_2311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_2312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_2313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_2314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_2315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_2316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_2317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_2318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_2319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_2320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_2321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_2322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_2323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_2324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_2325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_2326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_2327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_2328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_2329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_2330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_2331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_2332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_2333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_2334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_2335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_2336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_2337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_2339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_2340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_2343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_2346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_2347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_2348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_2349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_2350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_2351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_2352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_2353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_2354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_2355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_2356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_2357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_2358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_2359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_2360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_2361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_2362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_2363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_2364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_2365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_2366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_2367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_2368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_2369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_2370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_2371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_2372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_2374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_2375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_2378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_2381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_2382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_2383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_2384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_2385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_2386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_2387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_2388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_2389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_2390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_2391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_2392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_2393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_2394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_2395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_2396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_2397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_2398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_2399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_2400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_2401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_2402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_2403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_2404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_2405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_2406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_2407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_2408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_2410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_2411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_2412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_2414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_2417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_2418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_2419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_2420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_2421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_2422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_2423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_2424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_2425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_2426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_2427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_2428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_2429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_2430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_2431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_2432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_2433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_2434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_2435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_2436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_2437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_2438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_2439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_2440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_2441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_2442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_2443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_2445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_2446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_2447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_2449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_2450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_2452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_2453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_2454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_2455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_2456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_2457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_2458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_2459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_2460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_2461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_2462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_2463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_2464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_2465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_2466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_2467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_2468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_2469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_2470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_2471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_2472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_2473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_2474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_2475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_2476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_2477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_2478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_2479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_2481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_2482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_2483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_2485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_2486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_2488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_2489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_2490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_2491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_2492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_2493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_2494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_2495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_2497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_2498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_2499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_2500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_2501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_2502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_2503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_2504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_2505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_2506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_2507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_2508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_2509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_2510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_2511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_2512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_2513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_2514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_2516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_2517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_2518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_2520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_2521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_2523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_2524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_2525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_2526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_2529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_2530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_2531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_2532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_2533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_2534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_2535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_2536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_2537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_2539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_2540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_2541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_2542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_2543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_2544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_2545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_2546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_2547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_2548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_2549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_2550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_2552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_2553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_2556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_2560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_2561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_2563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_2564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_2565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_2566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_2567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_2568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_2569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_2570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_2571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_2572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_2573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_2574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_2575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_2576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_2577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_2578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_2579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_2580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_2581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_2582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_2583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_2584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_2585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_2587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_2588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_2594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_2596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_2597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_2599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_2600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_2601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_2602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_2603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_2604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_2605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_2606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_2607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_2608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_2609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_2610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_2611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_2612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_2613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_2614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_2615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_2616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_2617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_2618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_2619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_2620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_2623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_2624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_2627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_2628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_2631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_2632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_2634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_2635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_2636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_2637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_2638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_2639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_2640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_2643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_2644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_2646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_2647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_2648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_2650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_2652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_2653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_2654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_2655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_2656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_2658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_2659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_2660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_2663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_2665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_2667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_2668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_2670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_2671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_2672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_2673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_2674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_2675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_2676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_2677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_2678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_2679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_2680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_2681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_2682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_2683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_2684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_2686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_2687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_2688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_2689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_2690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_2691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_2692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_2694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_2695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_2696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_2698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_2701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_2702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_2703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_2704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_2705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_2706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_2707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_2708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_2709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_2710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_2711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_2712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_2713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_2714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_2715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_2716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_2717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_2718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_2719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_2720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_2721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_2722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_2723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_2724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_2725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_2726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_2727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_2729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_2730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_2731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_2733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_2734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_2736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_2737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_2738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_2739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_2740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_2741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_2742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_2743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_2744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_2745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_2746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_2747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_2748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_2749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_2750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_2751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_2752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_2753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_2754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_2755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_2756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_2757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_2758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_2759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_2760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_2761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_2762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_2763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_2765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_2766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_2767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_2769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_2770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_2772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_2773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_2774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_2775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_2776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_2777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_2778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_2779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_2780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_2781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_2782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_2783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_2784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_2785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_2786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_2787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_2788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_2789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_2790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_2791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_2792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_2793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_2794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_2795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_2796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_2797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_2798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_2800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_2801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_2802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_2804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_2805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_2807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_2808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_2809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_2810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_2811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_2812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_2813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_2814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_2816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_2817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_2818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_2819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_2820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_2821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_2822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_2823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_2824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_2825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_2826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_2827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_2828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_2829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_2830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_2831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_2832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_2833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_2834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_2836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_2837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_2838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_2840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_2843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_2844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_2845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_2846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_2849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_2851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_2852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_2853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_2854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_2856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_2858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_2859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_2860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_2861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_2862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_2863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_2864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_2865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_2866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_2867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_2868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_2869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_2871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_2872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_2873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_2875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_2876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_2878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_2879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_2881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_2882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_2884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_2885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_2886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_2887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_2888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_2889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_2890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_2891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_2892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_2893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_2894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_2895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_2896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_2897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_2898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_2899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_2900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_2901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_2902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_2903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_2904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_2905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_2907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_2908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_2909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_2911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_2914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_2915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_2917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_2918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_2920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_2921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_2922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_2923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_2924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_2925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_2926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_2927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_2928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_2929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_2930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_2931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_2932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_2933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_2934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_2935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_2936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_2937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_2938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_2939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_2940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_2942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_2943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_2944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_2946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_2949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_2950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_2952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_2953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_2955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_2956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_2957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_2958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_2959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_2960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_2961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_2962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_2963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_2964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_2965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_2966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_2967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_2968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_2969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_2970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_2971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_2972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_2973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_2974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_2975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_2976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_2978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_2979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_2980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_2982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_2985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_2988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_2989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_2991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_2992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_2993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_2994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_2995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_2996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_2997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_2998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_2999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_3000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_3001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_3003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_3004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_3005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_3007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_3009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_3010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_3011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_3013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_3014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_3015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_3017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_3018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_3020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_3021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_3022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_3023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_3024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_3025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_3026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_3028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_3029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_3030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_3031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_3032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_3033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_3034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_3035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_3036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_3037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_3038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_3039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_3040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_3041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_3042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_3043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_3044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_3045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_3046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_3047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_3049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_3050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_3051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_3053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_3054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_3056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_3057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_3058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_3060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_3061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_3063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_3064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_3065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_3066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_3067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_3068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_3069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_3070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_3071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_3072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_3073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_3074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_3075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_3076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_3077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_3078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_3079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_3080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_3081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_3082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_3084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_3085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_3086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_3088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_3089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_3092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_3093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_3094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_3096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_3097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_3099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_3100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_3101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_3102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_3103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_3104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_3105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_3106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_3107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_3108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_3109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_3110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_3111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_3112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_3113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_3114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_3115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_3116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_3117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_3118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_3120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_3121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_3122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_3124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_3125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_3127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_3128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_3129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_3131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_3132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_3135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_3136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_3137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_3138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_3139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_3140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_3141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_3142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_3143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_3144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_3145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_3146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_3147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_3148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_3149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_3150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_3151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_3152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_3153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_3155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_3156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_3157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_3159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_3160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_3163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_3164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_3165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_3167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_3168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_3170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_3171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_3172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_3176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_3178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_3179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_3180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_3181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_3183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_3184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_3188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_3189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_3190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_3191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_3192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_3194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_3195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_3196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_3198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_3200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_3201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_3202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_3203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_3204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_3205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_3206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_3207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_3208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_3209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_3210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_3211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_3212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_3213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_3214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_3215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_3216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_3217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_3218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_3219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_3220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_3221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_3222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_3223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_3224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_3225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_3226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_3227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_3228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_3229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_3230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_3231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_3232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_3233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_3234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_3235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_3236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_3237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_3238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_3239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_3240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_3241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_3242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_3243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_3244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_3245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_3246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_3247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_3248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_3249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_3250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_3251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_3252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_3253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_3254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_3255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_3256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_3257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_3258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_3259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_3260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_3261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_3262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_3263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_3264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_3265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_3266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_3267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_3268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_3269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_3270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_3271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_3272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_3273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_3274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_3275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_3276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_3277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_3278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_3279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_3280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_3281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_3282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_3283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_3284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_3285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_3286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_3287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_3288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_3289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_3290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_3291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_3292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_3293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_3294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_3295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_3296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_3297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_3298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_3299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_3300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_3301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_3302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_3303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_3304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_3305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_3306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_3307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_3308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_3309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_3310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_3311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_3312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_3313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_3314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_3315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_3316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_3317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_3318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_3319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_3320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_3321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_3322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_3323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_3324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_3325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_3326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_3327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_3328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_3329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_3330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_3331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_3332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_3333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_3334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_3335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_3336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_3337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_3338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_3339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_3340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_3341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_3342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_3343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_3344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_3345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_3346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_3347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_3348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_3349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_3350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_3351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_3352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_3353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_3354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_3355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_3356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_3357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_3358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_3359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_3360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_3361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_3362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_3363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_3364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_3365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_3366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_3367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_3368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_3369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_3370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_3371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_3372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_3373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_3374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_3375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_3376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_3377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_3378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_3379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_3380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_3381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_3382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_3383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_3384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_3385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_3386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_3387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_3388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_3389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_3390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_3391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_3392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_3393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_3394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_3395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_3396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_3397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_3398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_3399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_3400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_3401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_3402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_3403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_3404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_3405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_3406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_3407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_3408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_3409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_3410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_3411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_3412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_3413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_3414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_3415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_3416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_3417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_3418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_3419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_3420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_3421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_3422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_3423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_3424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_3425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_3426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_3427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_3428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_3429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_3430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_3431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_3432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_3433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_3434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_3435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_3436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_3437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_3438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_3439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_3440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_3441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_3442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_3443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_3444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_3445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_3446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_3447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_3448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_3449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_3450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_3451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_3452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_3454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_3455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_3456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_3457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_3458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_3459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_3460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_3461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_3462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_3463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_3464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_3465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_3466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_3467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_3468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_3469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_3470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_3471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_3472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_3473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_3474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_3475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_3476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_3477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_3478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_3479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_3480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_3481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_3482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_3483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_3484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_3486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_3487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_3489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_3490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_3491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_3493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_3495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_3496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_3497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_3498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_3499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_3500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_3501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_3502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_3503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_3504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_3505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_3506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_3507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_3508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_3509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_3510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_3511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_3512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_3513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_3514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_3515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_3516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_3517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_3518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_3519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_3520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_3521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_3522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_3523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_3524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_3525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_3526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_3527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_3528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_3529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_3530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_3531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_3532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_3533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_3534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_3535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_3536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_3537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_3538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_3539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_3540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_3541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_3542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_3543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_3544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_3545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_3546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_3547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_3548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_171_3549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_171_3550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_171_3551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_171_3552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_171_3553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_171_3554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_171_3555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_171_3556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_171_3557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_171_3558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_171_3559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_171_3560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_171_3561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_171_3562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_171_3563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_171_3564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_171_3565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_171_3566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_3567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_3568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_3569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_3570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_3571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_3572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_3573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_3574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_3575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_3576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_3577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_3578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_3579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_3580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_3581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_3582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_3583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_3584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_3585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_173_3586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_173_3587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_173_3588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_173_3589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_173_3590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_173_3591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_173_3592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_173_3593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_173_3594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_173_3595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_173_3596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_173_3597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_173_3598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_173_3599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_173_3600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_173_3601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_173_3602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_173_3603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_3604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_3605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_3606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_3607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_3608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_3609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_3610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_3611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_3612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_3613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_3614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_3615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_3616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_3617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_3618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_3619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_3620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_3621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_3622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_175_3623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_175_3624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_175_3625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_175_3626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_175_3627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_175_3628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_175_3629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_175_3630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_175_3631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_175_3632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_175_3633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_175_3634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_175_3635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_175_3636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_175_3637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_175_3638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_175_3639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_175_3640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_3641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_3642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_3643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_3644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_3645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_3646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_3647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_3648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_3649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_3650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_3651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_3652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_3653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_3654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_3655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_3656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_3657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_3658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_3659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_177_3660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_177_3661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_177_3662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_177_3663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_177_3664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_177_3665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_177_3666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_177_3667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_177_3668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_177_3669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_177_3670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_177_3671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_177_3672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_177_3673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_177_3674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_177_3675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_177_3676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_177_3677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_3678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_3679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_3680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_3681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_3682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_3683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_3684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_3685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_3686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_3687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_3688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_3689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_3690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_3691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_3692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_3693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_3694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_3695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_3696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_179_3697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_179_3698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_179_3699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_179_3700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_179_3701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_179_3702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_179_3703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_179_3704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_179_3705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_179_3706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_179_3707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_179_3708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_179_3709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_179_3710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_179_3711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_179_3712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_179_3713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_179_3714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_3715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_3716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_3717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_3718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_3719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_3720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_3721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_3722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_3723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_3724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_3725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_3726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_3727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_3728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_3729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_3730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_3731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_3732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_3733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_3734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_3735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_3736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_3737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_3738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_3739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_3740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_3741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_3742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_3743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_3744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_3745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_3746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_3747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_3748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_3749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_3750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_3751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_3752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_3753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_3754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_3755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_3756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_3757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_3758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_3759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_3760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_3761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_3762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_3763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_3764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_3765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_3766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_3767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_3768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_3769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_3770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_3772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_3773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_3774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_3775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_3776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_3777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_3778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_3779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_3780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_3781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_3782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_3783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_3784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_3785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_3786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_3787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_3788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_3789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_1958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_1959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_1960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_1961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_1962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_1963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_1964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_1965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_1966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_1967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_1968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_1969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_1970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_1971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_1972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_1973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_1974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_1975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_1995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_1996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_1997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_1998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_1999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_569 ();
 gf180mcu_fd_sc_mcu7t5v0__clkinv_3 _08467_ (.I(net4),
    .ZN(_00997_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _08468_ (.I(net5),
    .ZN(_00998_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _08469_ (.A1(net6),
    .A2(_00998_),
    .ZN(_00999_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _08470_ (.A1(_00997_),
    .A2(net3),
    .A3(_00999_),
    .ZN(_01000_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08471_ (.A1(net2),
    .A2(net1),
    .ZN(_01001_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08472_ (.A1(_01000_),
    .A2(_01001_),
    .ZN(_01002_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _08473_ (.A1(net7),
    .A2(net16),
    .Z(_01003_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08474_ (.A1(_01002_),
    .A2(_01003_),
    .Z(_01004_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08475_ (.I(_01004_),
    .Z(_01005_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _08476_ (.I(net13),
    .ZN(_01006_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08477_ (.A1(_01006_),
    .A2(_01005_),
    .ZN(_01007_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _08478_ (.A1(\filters.res_filt[5] ),
    .A2(_01005_),
    .B(_01007_),
    .ZN(_01008_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08479_ (.I(_01008_),
    .ZN(_01009_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08480_ (.I(net17),
    .Z(_01010_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08481_ (.A1(_01002_),
    .A2(_01003_),
    .ZN(_01011_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08482_ (.A1(net14),
    .A2(_01011_),
    .ZN(_01012_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08483_ (.I(_01004_),
    .Z(_01013_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08484_ (.A1(\filters.res_filt[6] ),
    .A2(_01013_),
    .ZN(_01014_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _08485_ (.A1(_01010_),
    .A2(_01012_),
    .A3(_01014_),
    .Z(_01015_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08486_ (.I(_01015_),
    .Z(_01016_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _08487_ (.I(net12),
    .ZN(_01017_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08488_ (.A1(_01017_),
    .A2(_01005_),
    .ZN(_01018_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _08489_ (.A1(\filters.res_filt[4] ),
    .A2(_01005_),
    .B(_01018_),
    .ZN(_01019_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08490_ (.A1(_01010_),
    .A2(_01019_),
    .ZN(_01020_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08491_ (.I(_01020_),
    .Z(_00129_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08492_ (.A1(_01016_),
    .A2(_00129_),
    .ZN(_01021_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08493_ (.A1(net15),
    .A2(_01011_),
    .ZN(_01022_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08494_ (.A1(\filters.res_filt[7] ),
    .A2(_01013_),
    .ZN(_01023_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _08495_ (.A1(_01010_),
    .A2(_01022_),
    .A3(_01023_),
    .Z(_01024_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08496_ (.I(_01024_),
    .Z(_01025_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08497_ (.I(_01015_),
    .ZN(_01026_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08498_ (.A1(_01026_),
    .A2(_01019_),
    .ZN(_01027_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08499_ (.A1(_01009_),
    .A2(_01021_),
    .B(_01025_),
    .C(_01027_),
    .ZN(_01028_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08500_ (.I(_01024_),
    .ZN(_01029_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08501_ (.I(_01029_),
    .Z(_00132_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08502_ (.I(_01026_),
    .Z(_01030_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08503_ (.A1(_01009_),
    .A2(_00129_),
    .ZN(_01031_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _08504_ (.I(_01010_),
    .Z(_01032_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _08505_ (.A1(_01008_),
    .A2(_01019_),
    .B(_01032_),
    .ZN(_01033_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08506_ (.A1(_01031_),
    .A2(_01033_),
    .ZN(_01034_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08507_ (.A1(_01030_),
    .A2(_01034_),
    .ZN(_01035_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08508_ (.I(_01031_),
    .Z(_01036_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08509_ (.A1(_01016_),
    .A2(_01036_),
    .ZN(_01037_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08510_ (.A1(_00132_),
    .A2(_01035_),
    .A3(_01037_),
    .ZN(_01038_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08511_ (.A1(_01028_),
    .A2(_01038_),
    .Z(_01039_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08512_ (.I(_01039_),
    .Z(_00000_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08513_ (.I(_01008_),
    .Z(_01040_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08514_ (.A1(_01040_),
    .A2(_01030_),
    .B(_00129_),
    .ZN(_01041_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _08515_ (.I(net17),
    .Z(_01042_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08516_ (.I(_01042_),
    .Z(_01043_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _08517_ (.A1(_01043_),
    .A2(_01008_),
    .B(_01016_),
    .ZN(_01044_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _08518_ (.A1(_01024_),
    .A2(_01027_),
    .A3(_01044_),
    .ZN(_01045_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08519_ (.A1(_01041_),
    .A2(_01045_),
    .Z(_01046_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08520_ (.I(_01046_),
    .Z(_00001_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08521_ (.A1(_01027_),
    .A2(_01036_),
    .B(_01029_),
    .ZN(_01047_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08522_ (.A1(_01021_),
    .A2(_01035_),
    .ZN(_01048_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08523_ (.I0(_01047_),
    .I1(_00132_),
    .S(_01048_),
    .Z(_01049_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08524_ (.I(_01049_),
    .Z(_00002_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08525_ (.I(_01025_),
    .Z(_01050_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08526_ (.A1(_01043_),
    .A2(_01040_),
    .ZN(_01051_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08527_ (.I(_01051_),
    .Z(_00130_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08528_ (.A1(_01027_),
    .A2(_01031_),
    .ZN(_01052_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08529_ (.A1(_01050_),
    .A2(_00130_),
    .B(_01052_),
    .ZN(_01053_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08530_ (.A1(_01047_),
    .A2(_01053_),
    .Z(_01054_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08531_ (.I(_01054_),
    .Z(_00003_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08532_ (.A1(_01016_),
    .A2(_00130_),
    .ZN(_01055_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08533_ (.A1(_01040_),
    .A2(_01030_),
    .B(_01025_),
    .ZN(_01056_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08534_ (.A1(_01021_),
    .A2(_01055_),
    .A3(_01056_),
    .ZN(_01057_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08535_ (.I(_01030_),
    .Z(_00131_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08536_ (.A1(_00131_),
    .A2(_01050_),
    .A3(_01036_),
    .ZN(_01058_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08537_ (.A1(_01057_),
    .A2(_01058_),
    .ZN(_00004_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08538_ (.A1(_01036_),
    .A2(_01044_),
    .ZN(_01059_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08539_ (.I0(_01019_),
    .I1(_01059_),
    .S(_01025_),
    .Z(_01060_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08540_ (.I(_01060_),
    .Z(_00005_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08541_ (.A1(_01040_),
    .A2(_01050_),
    .B(_01045_),
    .ZN(_00006_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08542_ (.A1(_01050_),
    .A2(_01048_),
    .B1(_01055_),
    .B2(_01056_),
    .ZN(_00007_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08543_ (.A1(_00131_),
    .A2(_01033_),
    .ZN(_01061_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08544_ (.A1(_00132_),
    .A2(_01061_),
    .B(_01044_),
    .ZN(_00008_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _08545_ (.I(net17),
    .ZN(_01062_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08546_ (.I(\clk_ctr[0] ),
    .ZN(_01063_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _08547_ (.A1(\clk_trg[0] ),
    .A2(_01063_),
    .B(\clk_ctr[1] ),
    .ZN(_01064_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08548_ (.I(\clk_trg[1] ),
    .ZN(_01065_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08549_ (.A1(_01065_),
    .A2(\clk_ctr[1] ),
    .ZN(_01066_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08550_ (.A1(\clk_ctr[0] ),
    .A2(_01066_),
    .ZN(_01067_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _08551_ (.A1(\clk_trg[1] ),
    .A2(_01064_),
    .B1(_01067_),
    .B2(\clk_trg[0] ),
    .ZN(_01068_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _08552_ (.A1(_01062_),
    .A2(_01068_),
    .ZN(_01069_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08553_ (.A1(\channels.clk_div[0] ),
    .A2(_01069_),
    .ZN(_01070_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08554_ (.I(\channels.clk_div[2] ),
    .ZN(_01071_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08555_ (.I(\channels.clk_div[1] ),
    .Z(_01072_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08556_ (.A1(_01071_),
    .A2(_01072_),
    .ZN(_01073_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08557_ (.I(_01073_),
    .Z(_01074_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08558_ (.I(_01074_),
    .Z(_01075_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08559_ (.I(_01075_),
    .Z(_01076_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08560_ (.I(_01076_),
    .Z(_01077_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08561_ (.I(_01077_),
    .Z(_01078_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08562_ (.I(_01078_),
    .Z(_01079_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08563_ (.I(_01079_),
    .Z(_01080_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08564_ (.I(_01080_),
    .Z(_01081_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08565_ (.I(_01081_),
    .Z(_01082_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08566_ (.A1(_01070_),
    .A2(_01082_),
    .Z(_01083_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08567_ (.I(_01083_),
    .Z(_01084_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _08568_ (.I0(\channels.accum[0][23] ),
    .I1(\channels.accum[1][23] ),
    .I2(\channels.accum[2][23] ),
    .I3(\channels.accum[3][23] ),
    .S0(_00009_),
    .S1(_00010_),
    .Z(_01085_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08569_ (.I(_01085_),
    .Z(_01086_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08570_ (.I(_01042_),
    .Z(_01087_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08571_ (.A1(_01087_),
    .A2(_01083_),
    .ZN(_01088_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08572_ (.I(_01088_),
    .Z(_01089_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08573_ (.I(_01089_),
    .Z(_01090_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08574_ (.A1(_01084_),
    .A2(_01086_),
    .B1(_01090_),
    .B2(\channels.ring_outs[2] ),
    .ZN(_01091_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08575_ (.I(_01091_),
    .ZN(_00011_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _08576_ (.I(\channels.clk_div[0] ),
    .ZN(_01092_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _08577_ (.I(_01068_),
    .ZN(_01093_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08578_ (.A1(net17),
    .A2(_01093_),
    .ZN(_01094_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08579_ (.A1(_01092_),
    .A2(_01094_),
    .ZN(_01095_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08580_ (.I(_01071_),
    .Z(_01096_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08581_ (.I(_01096_),
    .Z(_01097_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08582_ (.I(_01072_),
    .Z(_01098_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08583_ (.A1(_01097_),
    .A2(_01098_),
    .ZN(_01099_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08584_ (.A1(_01095_),
    .A2(_01099_),
    .ZN(_01100_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08585_ (.I(_01100_),
    .Z(_01101_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08586_ (.I(_01042_),
    .Z(_01102_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08587_ (.A1(_01102_),
    .A2(_01100_),
    .ZN(_01103_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08588_ (.I(_01103_),
    .Z(_01104_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08589_ (.I(_01104_),
    .Z(_01105_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08590_ (.A1(_01086_),
    .A2(_01101_),
    .B1(_01105_),
    .B2(\channels.ring_outs[1] ),
    .ZN(_01106_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08591_ (.I(_01106_),
    .ZN(_00012_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08592_ (.I(\channels.lfsr[3][0] ),
    .Z(_01107_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08593_ (.I(_01107_),
    .Z(_00013_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08594_ (.I(\channels.lfsr[3][1] ),
    .Z(_01108_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08595_ (.I(_01108_),
    .Z(_00014_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08596_ (.I(\channels.lfsr[3][2] ),
    .Z(_01109_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08597_ (.I(_01109_),
    .Z(_00015_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08598_ (.I(\channels.lfsr[3][3] ),
    .Z(_01110_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08599_ (.I(_01110_),
    .Z(_00016_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08600_ (.I(\channels.lfsr[3][4] ),
    .Z(_01111_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08601_ (.I(_01111_),
    .Z(_00017_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08602_ (.I(\channels.lfsr[3][5] ),
    .Z(_01112_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08603_ (.I(_01112_),
    .Z(_00018_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08604_ (.I(\channels.lfsr[3][6] ),
    .Z(_01113_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08605_ (.I(_01113_),
    .Z(_00019_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08606_ (.I(\channels.lfsr[3][7] ),
    .Z(_01114_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08607_ (.I(_01114_),
    .Z(_00020_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08608_ (.I(\channels.lfsr[3][8] ),
    .Z(_01115_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08609_ (.I(_01115_),
    .Z(_00021_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08610_ (.I(\channels.lfsr[3][9] ),
    .Z(_01116_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08611_ (.I(_01116_),
    .Z(_00022_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08612_ (.I(\channels.lfsr[3][10] ),
    .Z(_01117_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08613_ (.I(_01117_),
    .Z(_00023_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08614_ (.I(\channels.lfsr[3][11] ),
    .Z(_01118_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08615_ (.I(_01118_),
    .Z(_00024_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08616_ (.I(\channels.lfsr[3][12] ),
    .Z(_01119_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08617_ (.I(_01119_),
    .Z(_00025_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08618_ (.I(\channels.lfsr[3][13] ),
    .Z(_01120_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08619_ (.I(_01120_),
    .Z(_00026_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08620_ (.I(\channels.lfsr[3][14] ),
    .Z(_01121_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08621_ (.I(_01121_),
    .Z(_00027_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08622_ (.I(\channels.lfsr[3][15] ),
    .Z(_01122_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08623_ (.I(_01122_),
    .Z(_00028_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08624_ (.I(\channels.lfsr[3][16] ),
    .Z(_01123_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08625_ (.I(_01123_),
    .Z(_00029_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08626_ (.I(\channels.lfsr[3][17] ),
    .Z(_01124_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08627_ (.I(_01124_),
    .Z(_00030_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08628_ (.I(\channels.lfsr[3][18] ),
    .Z(_01125_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08629_ (.I(_01125_),
    .Z(_00031_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08630_ (.I(\channels.lfsr[3][19] ),
    .Z(_01126_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08631_ (.I(_01126_),
    .Z(_00032_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08632_ (.I(\channels.lfsr[3][20] ),
    .Z(_01127_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08633_ (.I(_01127_),
    .Z(_00033_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08634_ (.I(\channels.lfsr[3][21] ),
    .Z(_01128_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08635_ (.I(_01128_),
    .Z(_00034_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08636_ (.I(\channels.lfsr[3][22] ),
    .Z(_01129_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08637_ (.I(_01129_),
    .Z(_00035_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08638_ (.I(\channels.env_vol[3][0] ),
    .Z(_01130_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08639_ (.I(_01130_),
    .Z(_00036_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08640_ (.I(\channels.env_vol[3][1] ),
    .Z(_01131_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08641_ (.I(_01131_),
    .Z(_00037_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08642_ (.I(\channels.env_vol[3][2] ),
    .Z(_01132_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08643_ (.I(_01132_),
    .Z(_00038_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08644_ (.I(\channels.env_vol[3][3] ),
    .Z(_01133_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08645_ (.I(_01133_),
    .Z(_00039_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08646_ (.I(\channels.env_vol[3][4] ),
    .Z(_01134_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08647_ (.I(_01134_),
    .Z(_00040_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08648_ (.I(\channels.env_vol[3][5] ),
    .Z(_01135_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08649_ (.I(_01135_),
    .Z(_00041_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08650_ (.I(\channels.env_vol[3][6] ),
    .Z(_01136_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08651_ (.I(_01136_),
    .Z(_00042_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08652_ (.I(\channels.env_vol[3][7] ),
    .Z(_01137_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08653_ (.I(_01137_),
    .Z(_00043_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08654_ (.I(_00009_),
    .Z(_01138_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08655_ (.I(_01138_),
    .Z(_01139_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _08656_ (.I(_01139_),
    .Z(_01140_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08657_ (.I(_01140_),
    .Z(_01141_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08658_ (.I(_01141_),
    .Z(_01142_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08659_ (.I(_01142_),
    .Z(_01143_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08660_ (.I(_01143_),
    .Z(_01144_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08661_ (.I(_01144_),
    .Z(_01145_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08662_ (.I(_01145_),
    .Z(_01146_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _08663_ (.I(_01146_),
    .Z(_01147_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08664_ (.I(_01147_),
    .Z(_01148_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08665_ (.I(_01148_),
    .Z(_01149_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08666_ (.I(_01149_),
    .Z(_01150_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08667_ (.I(_01150_),
    .Z(_01151_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _08668_ (.I(_01151_),
    .Z(_01152_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08669_ (.I(_00010_),
    .Z(_01153_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08670_ (.I(_01153_),
    .Z(_01154_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08671_ (.I(_01154_),
    .Z(_01155_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08672_ (.I(_01155_),
    .Z(_01156_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08673_ (.I(_01156_),
    .Z(_01157_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08674_ (.I(_01157_),
    .Z(_01158_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08675_ (.I(_01158_),
    .Z(_01159_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08676_ (.I(_01159_),
    .Z(_01160_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08677_ (.I(_01160_),
    .Z(_01161_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08678_ (.I(_01161_),
    .Z(_01162_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08679_ (.I(_01162_),
    .Z(_01163_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _08680_ (.I(_01163_),
    .Z(_01164_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08681_ (.I(_01164_),
    .Z(_01165_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08682_ (.I(_01165_),
    .Z(_01166_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08683_ (.I(_01166_),
    .Z(_01167_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _08684_ (.I(_01167_),
    .Z(_01168_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _08685_ (.I0(\channels.exp_counter[0][0] ),
    .I1(\channels.exp_counter[1][0] ),
    .I2(\channels.exp_counter[2][0] ),
    .I3(\channels.exp_counter[3][0] ),
    .S0(_01152_),
    .S1(_01168_),
    .Z(_01169_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08686_ (.I(_01165_),
    .Z(_01170_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08687_ (.I(_01170_),
    .Z(_01171_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08688_ (.I(_01171_),
    .Z(_01172_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08689_ (.I(_01172_),
    .Z(_01173_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08690_ (.I(_01173_),
    .Z(_01174_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08691_ (.I(_01152_),
    .Z(_01175_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08692_ (.I(_01175_),
    .Z(_01176_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08693_ (.I0(\channels.exp_periods[0][0] ),
    .I1(\channels.exp_periods[1][0] ),
    .S(_01176_),
    .Z(_01177_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08694_ (.I(_01175_),
    .Z(_01178_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08695_ (.I(_01178_),
    .Z(_01179_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08696_ (.I(\channels.exp_periods[2][0] ),
    .ZN(_01180_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08697_ (.A1(_01176_),
    .A2(\channels.exp_periods[3][0] ),
    .ZN(_01181_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _08698_ (.A1(_01179_),
    .A2(_01180_),
    .B(_01181_),
    .C(_01173_),
    .ZN(_01182_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _08699_ (.A1(_01174_),
    .A2(_01177_),
    .B(_01182_),
    .ZN(_01183_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08700_ (.A1(_01169_),
    .A2(_01183_),
    .ZN(_01184_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _08701_ (.I0(\channels.exp_counter[0][2] ),
    .I1(\channels.exp_counter[1][2] ),
    .I2(\channels.exp_counter[2][2] ),
    .I3(\channels.exp_counter[3][2] ),
    .S0(_01175_),
    .S1(_01172_),
    .Z(_01185_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08702_ (.I(_01185_),
    .Z(_01186_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08703_ (.I(_01178_),
    .Z(_01187_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08704_ (.I(_01173_),
    .Z(_01188_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _08705_ (.I0(\channels.exp_periods[0][2] ),
    .I1(\channels.exp_periods[1][2] ),
    .I2(\channels.exp_periods[2][2] ),
    .I3(\channels.exp_periods[3][2] ),
    .S0(_01187_),
    .S1(_01188_),
    .Z(_01189_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08706_ (.A1(_01186_),
    .A2(_01189_),
    .Z(_01190_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _08707_ (.I0(\channels.exp_counter[0][4] ),
    .I1(\channels.exp_counter[1][4] ),
    .I2(\channels.exp_counter[2][4] ),
    .I3(\channels.exp_counter[3][4] ),
    .S0(_01175_),
    .S1(_01172_),
    .Z(_01191_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08708_ (.I0(\channels.exp_periods[0][4] ),
    .I1(\channels.exp_periods[1][4] ),
    .S(_01178_),
    .Z(_01192_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08709_ (.I(\channels.exp_periods[2][4] ),
    .ZN(_01193_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08710_ (.A1(_01176_),
    .A2(\channels.exp_periods[3][4] ),
    .ZN(_01194_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _08711_ (.A1(_01179_),
    .A2(_01193_),
    .B(_01194_),
    .C(_01173_),
    .ZN(_01195_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _08712_ (.A1(_01174_),
    .A2(_01192_),
    .B(_01195_),
    .ZN(_01196_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08713_ (.A1(_01191_),
    .A2(_01196_),
    .Z(_01197_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _08714_ (.I0(\channels.exp_counter[0][3] ),
    .I1(\channels.exp_counter[1][3] ),
    .I2(\channels.exp_counter[2][3] ),
    .I3(\channels.exp_counter[3][3] ),
    .S0(_01178_),
    .S1(_01172_),
    .Z(_01198_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08715_ (.I(_01198_),
    .Z(_01199_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08716_ (.I0(\channels.exp_periods[0][3] ),
    .I1(\channels.exp_periods[1][3] ),
    .S(_01187_),
    .Z(_01200_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08717_ (.I(_01176_),
    .Z(_01201_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08718_ (.I(\channels.exp_periods[2][3] ),
    .ZN(_01202_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08719_ (.A1(_01179_),
    .A2(\channels.exp_periods[3][3] ),
    .ZN(_01203_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _08720_ (.A1(_01201_),
    .A2(_01202_),
    .B(_01203_),
    .C(_01188_),
    .ZN(_01204_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _08721_ (.A1(_01174_),
    .A2(_01200_),
    .B(_01204_),
    .ZN(_01205_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _08722_ (.I0(\channels.exp_counter[0][1] ),
    .I1(\channels.exp_counter[1][1] ),
    .I2(\channels.exp_counter[2][1] ),
    .I3(\channels.exp_counter[3][1] ),
    .S0(_01152_),
    .S1(_01168_),
    .Z(_01206_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08723_ (.I0(\channels.exp_periods[0][1] ),
    .I1(\channels.exp_periods[1][1] ),
    .S(_01187_),
    .Z(_01207_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08724_ (.I(\channels.exp_periods[2][1] ),
    .ZN(_01208_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08725_ (.A1(_01187_),
    .A2(\channels.exp_periods[3][1] ),
    .ZN(_01209_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _08726_ (.A1(_01179_),
    .A2(_01208_),
    .B(_01209_),
    .C(_01188_),
    .ZN(_01210_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _08727_ (.A1(_01174_),
    .A2(_01207_),
    .B(_01210_),
    .ZN(_01211_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08728_ (.A1(_01199_),
    .A2(_01205_),
    .B1(_01206_),
    .B2(_01211_),
    .ZN(_01212_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _08729_ (.A1(_01199_),
    .A2(_01205_),
    .B1(_01206_),
    .B2(_01211_),
    .ZN(_01213_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08730_ (.I(_01213_),
    .ZN(_01214_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08731_ (.A1(_01197_),
    .A2(_01212_),
    .A3(_01214_),
    .ZN(_01215_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _08732_ (.A1(_01184_),
    .A2(_01190_),
    .A3(_01215_),
    .ZN(_01216_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08733_ (.I(_01216_),
    .Z(_01217_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08734_ (.A1(_01169_),
    .A2(_01217_),
    .ZN(_01218_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08735_ (.I(_01100_),
    .Z(_01219_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08736_ (.I(_01219_),
    .Z(_01220_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08737_ (.A1(\channels.exp_counter[1][0] ),
    .A2(_01105_),
    .B1(_01218_),
    .B2(_01220_),
    .ZN(_01221_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08738_ (.I(_01221_),
    .ZN(_00044_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08739_ (.A1(_01169_),
    .A2(_01206_),
    .ZN(_01222_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08740_ (.A1(_01169_),
    .A2(_01206_),
    .Z(_01223_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08741_ (.A1(_01222_),
    .A2(_01223_),
    .ZN(_01224_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08742_ (.A1(_01217_),
    .A2(_01224_),
    .ZN(_01225_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08743_ (.A1(\channels.exp_counter[1][1] ),
    .A2(_01105_),
    .B1(_01225_),
    .B2(_01220_),
    .ZN(_01226_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08744_ (.I(_01226_),
    .ZN(_00045_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08745_ (.A1(_01186_),
    .A2(_01222_),
    .Z(_01227_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08746_ (.A1(_01217_),
    .A2(_01227_),
    .ZN(_01228_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08747_ (.A1(\channels.exp_counter[1][2] ),
    .A2(_01105_),
    .B1(_01228_),
    .B2(_01220_),
    .ZN(_01229_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08748_ (.I(_01229_),
    .ZN(_00046_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08749_ (.I(_01103_),
    .Z(_01230_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08750_ (.I(_01222_),
    .ZN(_01231_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08751_ (.A1(_01186_),
    .A2(_01199_),
    .A3(_01231_),
    .ZN(_01232_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08752_ (.A1(_01186_),
    .A2(_01231_),
    .B(_01199_),
    .ZN(_01233_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08753_ (.A1(_01216_),
    .A2(_01233_),
    .ZN(_01234_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08754_ (.A1(_01232_),
    .A2(_01234_),
    .Z(_01235_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08755_ (.A1(\channels.exp_counter[1][3] ),
    .A2(_01230_),
    .B1(_01235_),
    .B2(_01220_),
    .ZN(_01236_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08756_ (.I(_01236_),
    .ZN(_00047_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08757_ (.A1(_01191_),
    .A2(_01232_),
    .Z(_01237_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08758_ (.A1(_01217_),
    .A2(_01237_),
    .ZN(_01238_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08759_ (.A1(\channels.exp_counter[1][4] ),
    .A2(_01230_),
    .B1(_01238_),
    .B2(_01101_),
    .ZN(_01239_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08760_ (.I(_01239_),
    .ZN(_00048_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08761_ (.I(_01083_),
    .Z(_01240_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08762_ (.I(_01240_),
    .Z(_01241_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08763_ (.A1(\channels.exp_counter[2][0] ),
    .A2(_01090_),
    .B1(_01218_),
    .B2(_01241_),
    .ZN(_01242_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08764_ (.I(_01242_),
    .ZN(_00049_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08765_ (.A1(\channels.exp_counter[2][1] ),
    .A2(_01090_),
    .B1(_01225_),
    .B2(_01241_),
    .ZN(_01243_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08766_ (.I(_01243_),
    .ZN(_00050_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08767_ (.A1(\channels.exp_counter[2][2] ),
    .A2(_01090_),
    .B1(_01228_),
    .B2(_01241_),
    .ZN(_01244_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08768_ (.I(_01244_),
    .ZN(_00051_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08769_ (.I(_01088_),
    .Z(_01245_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08770_ (.A1(\channels.exp_counter[2][3] ),
    .A2(_01245_),
    .B1(_01235_),
    .B2(_01241_),
    .ZN(_01246_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08771_ (.I(_01246_),
    .ZN(_00052_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08772_ (.A1(\channels.exp_counter[2][4] ),
    .A2(_01245_),
    .B1(_01238_),
    .B2(_01084_),
    .ZN(_01247_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08773_ (.I(_01247_),
    .ZN(_00053_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08774_ (.I(\channels.clk_div[2] ),
    .Z(_01248_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08775_ (.I(_01248_),
    .Z(_01249_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08776_ (.I(_01072_),
    .Z(_01250_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08777_ (.A1(_01249_),
    .A2(_01250_),
    .Z(_01251_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08778_ (.I(_01251_),
    .Z(_01252_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08779_ (.A1(_01095_),
    .A2(_01252_),
    .ZN(_01253_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08780_ (.I(_01253_),
    .Z(_01254_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08781_ (.I(_01254_),
    .Z(_01255_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08782_ (.A1(_01102_),
    .A2(_01253_),
    .ZN(_01256_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08783_ (.I(_01256_),
    .Z(_01257_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08784_ (.I(_01257_),
    .Z(_01258_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08785_ (.A1(_01086_),
    .A2(_01255_),
    .B1(_01258_),
    .B2(\channels.ring_outs[0] ),
    .ZN(_01259_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08786_ (.I(_01259_),
    .ZN(_00054_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08787_ (.I(\channels.accum[0][0] ),
    .ZN(_01260_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08788_ (.I(_01256_),
    .Z(_01261_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08789_ (.I(_01261_),
    .Z(_01262_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08790_ (.I(_01250_),
    .Z(_01263_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _08791_ (.I(_01263_),
    .Z(_01264_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08792_ (.I(_01096_),
    .Z(_01265_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08793_ (.I(_01265_),
    .Z(_01266_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08794_ (.I(_01266_),
    .Z(_01267_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08795_ (.A1(_01267_),
    .A2(\channels.ctrl_reg2[3] ),
    .ZN(_01268_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _08796_ (.A1(_01267_),
    .A2(\channels.ctrl_reg3[3] ),
    .B1(\channels.ctrl_reg1[3] ),
    .B2(_01252_),
    .ZN(_01269_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _08797_ (.A1(_01264_),
    .A2(_01268_),
    .B(_01269_),
    .ZN(_01270_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08798_ (.A1(\channels.ctrl_reg3[1] ),
    .A2(\channels.sync_outs[1] ),
    .A3(_01082_),
    .ZN(_01271_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _08799_ (.I(\channels.clk_div[1] ),
    .ZN(_01272_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08800_ (.A1(_01248_),
    .A2(_01272_),
    .ZN(_01273_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08801_ (.I(_01273_),
    .Z(_01274_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08802_ (.I(_01274_),
    .Z(_01275_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08803_ (.I(_01275_),
    .Z(_01276_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08804_ (.I(_01276_),
    .Z(_01277_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08805_ (.I(_01277_),
    .Z(_01278_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08806_ (.I(_01278_),
    .Z(_01279_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08807_ (.I(_01279_),
    .Z(_01280_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _08808_ (.I(_01280_),
    .Z(_01281_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08809_ (.I(_01281_),
    .Z(_01282_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08810_ (.A1(\channels.ctrl_reg2[1] ),
    .A2(\channels.sync_outs[0] ),
    .A3(_01282_),
    .ZN(_01283_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08811_ (.A1(_01248_),
    .A2(\channels.clk_div[1] ),
    .ZN(_01284_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08812_ (.I(_01284_),
    .Z(_01285_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08813_ (.I(_01285_),
    .Z(_01286_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08814_ (.I(_01286_),
    .Z(_01287_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08815_ (.I(_01287_),
    .Z(_01288_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08816_ (.I(_01288_),
    .Z(_01289_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08817_ (.I(_01289_),
    .Z(_01290_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08818_ (.I(_01290_),
    .Z(_01291_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08819_ (.I(_01291_),
    .Z(_01292_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08820_ (.I(_01292_),
    .Z(_01293_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08821_ (.I(_01293_),
    .Z(_01294_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08822_ (.I(_01294_),
    .Z(_01295_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08823_ (.A1(\channels.ctrl_reg1[1] ),
    .A2(\channels.sync_outs[2] ),
    .A3(_01295_),
    .ZN(_01296_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08824_ (.A1(_01271_),
    .A2(_01283_),
    .A3(_01296_),
    .ZN(_01297_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08825_ (.A1(_01270_),
    .A2(_01297_),
    .ZN(_01298_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08826_ (.I(_01298_),
    .Z(_01299_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08827_ (.I(_01299_),
    .Z(_01300_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08828_ (.A1(\channels.freq3[0] ),
    .A2(_01074_),
    .ZN(_01301_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _08829_ (.A1(\channels.freq2[0] ),
    .A2(_01274_),
    .B1(_01287_),
    .B2(\channels.freq1[0] ),
    .ZN(_01302_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08830_ (.A1(_01301_),
    .A2(_01302_),
    .ZN(_01303_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08831_ (.I(_01188_),
    .Z(_01304_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08832_ (.I(_01142_),
    .Z(_01305_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08833_ (.I(_01305_),
    .Z(_01306_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08834_ (.I(_01306_),
    .Z(_01307_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08835_ (.I(_01307_),
    .Z(_01308_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08836_ (.A1(_01308_),
    .A2(\channels.accum[1][0] ),
    .ZN(_01309_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08837_ (.A1(_01146_),
    .A2(_01260_),
    .B(_01309_),
    .ZN(_01310_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08838_ (.I(\channels.accum[2][0] ),
    .ZN(_01311_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08839_ (.A1(_01308_),
    .A2(\channels.accum[3][0] ),
    .ZN(_01312_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _08840_ (.A1(_01308_),
    .A2(_01311_),
    .B(_01312_),
    .C(_01159_),
    .ZN(_01313_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08841_ (.A1(_01304_),
    .A2(_01310_),
    .B(_01313_),
    .ZN(_01314_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08842_ (.A1(_01303_),
    .A2(_01314_),
    .ZN(_01315_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08843_ (.A1(_01300_),
    .A2(_01315_),
    .ZN(_01316_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08844_ (.I(_01253_),
    .Z(_01317_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08845_ (.I(_01317_),
    .Z(_01318_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08846_ (.A1(_01260_),
    .A2(_01262_),
    .B1(_01316_),
    .B2(_01318_),
    .ZN(_00055_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08847_ (.I(_01295_),
    .Z(_01319_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08848_ (.A1(_01070_),
    .A2(_01319_),
    .ZN(_01320_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08849_ (.I(_01320_),
    .Z(_01321_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08850_ (.I(_01321_),
    .Z(_01322_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08851_ (.I(_01298_),
    .Z(_01323_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08852_ (.A1(_01160_),
    .A2(_01310_),
    .B(_01313_),
    .C(_01303_),
    .ZN(_01324_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08853_ (.A1(\channels.freq3[1] ),
    .A2(_01074_),
    .ZN(_01325_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _08854_ (.A1(\channels.freq2[1] ),
    .A2(_01274_),
    .B1(_01287_),
    .B2(\channels.freq1[1] ),
    .ZN(_01326_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08855_ (.A1(_01325_),
    .A2(_01326_),
    .ZN(_01327_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08856_ (.I(_01158_),
    .Z(_01328_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _08857_ (.I0(\channels.accum[0][1] ),
    .I1(\channels.accum[1][1] ),
    .I2(\channels.accum[2][1] ),
    .I3(\channels.accum[3][1] ),
    .S0(_01307_),
    .S1(_01328_),
    .Z(_01329_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08858_ (.A1(_01327_),
    .A2(_01329_),
    .ZN(_01330_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08859_ (.A1(_01324_),
    .A2(_01330_),
    .ZN(_01331_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08860_ (.A1(_01324_),
    .A2(_01330_),
    .Z(_01332_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _08861_ (.A1(_01323_),
    .A2(_01331_),
    .A3(_01332_),
    .ZN(_01333_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08862_ (.I(_01256_),
    .Z(_01334_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08863_ (.A1(\channels.accum[0][1] ),
    .A2(_01334_),
    .ZN(_01335_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08864_ (.A1(_01322_),
    .A2(_01333_),
    .B(_01335_),
    .ZN(_00056_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08865_ (.I(\channels.accum[0][2] ),
    .ZN(_01336_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08866_ (.I(_01299_),
    .Z(_01337_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08867_ (.A1(_01327_),
    .A2(_01329_),
    .ZN(_01338_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08868_ (.A1(\channels.freq3[2] ),
    .A2(_01075_),
    .ZN(_01339_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _08869_ (.A1(\channels.freq2[2] ),
    .A2(_01275_),
    .B1(_01287_),
    .B2(\channels.freq1[2] ),
    .ZN(_01340_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08870_ (.A1(_01339_),
    .A2(_01340_),
    .ZN(_01341_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _08871_ (.I0(\channels.accum[0][2] ),
    .I1(\channels.accum[1][2] ),
    .I2(\channels.accum[2][2] ),
    .I3(\channels.accum[3][2] ),
    .S0(_01145_),
    .S1(_01159_),
    .Z(_01342_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08872_ (.A1(_01341_),
    .A2(_01342_),
    .ZN(_01343_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08873_ (.A1(_01338_),
    .A2(_01332_),
    .A3(_01343_),
    .ZN(_01344_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08874_ (.A1(_01338_),
    .A2(_01332_),
    .ZN(_01345_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08875_ (.I(_01343_),
    .ZN(_01346_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08876_ (.A1(_01345_),
    .A2(_01346_),
    .ZN(_01347_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _08877_ (.A1(_01337_),
    .A2(_01344_),
    .A3(_01347_),
    .ZN(_01348_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08878_ (.A1(_01336_),
    .A2(_01262_),
    .B1(_01348_),
    .B2(_01318_),
    .ZN(_00057_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08879_ (.I(_01299_),
    .Z(_01349_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08880_ (.A1(_01341_),
    .A2(_01342_),
    .ZN(_01350_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08881_ (.A1(_01350_),
    .A2(_01347_),
    .ZN(_01351_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08882_ (.A1(\channels.freq3[3] ),
    .A2(_01075_),
    .ZN(_01352_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _08883_ (.A1(\channels.freq2[3] ),
    .A2(_01275_),
    .B1(_01288_),
    .B2(\channels.freq1[3] ),
    .ZN(_01353_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08884_ (.A1(_01352_),
    .A2(_01353_),
    .ZN(_01354_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _08885_ (.I0(\channels.accum[0][3] ),
    .I1(\channels.accum[1][3] ),
    .I2(\channels.accum[2][3] ),
    .I3(\channels.accum[3][3] ),
    .S0(_01308_),
    .S1(_01160_),
    .Z(_01355_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08886_ (.A1(_01354_),
    .A2(_01355_),
    .ZN(_01356_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08887_ (.I(_01356_),
    .ZN(_01357_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08888_ (.A1(_01351_),
    .A2(_01357_),
    .Z(_01358_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08889_ (.A1(_01349_),
    .A2(_01358_),
    .ZN(_01359_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08890_ (.I(_01257_),
    .Z(_01360_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08891_ (.A1(\channels.accum[0][3] ),
    .A2(_01360_),
    .ZN(_01361_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08892_ (.A1(_01322_),
    .A2(_01359_),
    .B(_01361_),
    .ZN(_00058_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08893_ (.I(\channels.accum[0][4] ),
    .ZN(_01362_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08894_ (.A1(_01350_),
    .A2(_01347_),
    .B(_01356_),
    .ZN(_01363_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08895_ (.A1(_01354_),
    .A2(_01355_),
    .B(_01363_),
    .ZN(_01364_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08896_ (.A1(\channels.freq3[4] ),
    .A2(_01075_),
    .ZN(_01365_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _08897_ (.A1(\channels.freq2[4] ),
    .A2(_01275_),
    .B1(_01288_),
    .B2(\channels.freq1[4] ),
    .ZN(_01366_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08898_ (.A1(_01365_),
    .A2(_01366_),
    .ZN(_01367_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _08899_ (.I0(\channels.accum[0][4] ),
    .I1(\channels.accum[1][4] ),
    .I2(\channels.accum[2][4] ),
    .I3(\channels.accum[3][4] ),
    .S0(_01146_),
    .S1(_01161_),
    .Z(_01368_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08900_ (.A1(_01367_),
    .A2(_01368_),
    .ZN(_01369_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08901_ (.A1(_01364_),
    .A2(_01369_),
    .ZN(_01370_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08902_ (.A1(_01364_),
    .A2(_01369_),
    .Z(_01371_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _08903_ (.A1(_01337_),
    .A2(_01370_),
    .A3(_01371_),
    .ZN(_01372_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08904_ (.A1(_01362_),
    .A2(_01262_),
    .B1(_01372_),
    .B2(_01318_),
    .ZN(_00059_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08905_ (.A1(_01367_),
    .A2(_01368_),
    .ZN(_01373_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08906_ (.A1(_01373_),
    .A2(_01371_),
    .ZN(_01374_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08907_ (.A1(\channels.freq3[5] ),
    .A2(_01076_),
    .ZN(_01375_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _08908_ (.A1(\channels.freq2[5] ),
    .A2(_01276_),
    .B1(_01288_),
    .B2(\channels.freq1[5] ),
    .ZN(_01376_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08909_ (.A1(_01375_),
    .A2(_01376_),
    .ZN(_01377_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _08910_ (.I0(\channels.accum[0][5] ),
    .I1(\channels.accum[1][5] ),
    .I2(\channels.accum[2][5] ),
    .I3(\channels.accum[3][5] ),
    .S0(_01147_),
    .S1(_01161_),
    .Z(_01378_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08911_ (.A1(_01377_),
    .A2(_01378_),
    .ZN(_01379_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08912_ (.A1(_01374_),
    .A2(_01379_),
    .ZN(_01380_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08913_ (.A1(_01349_),
    .A2(_01380_),
    .ZN(_01381_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08914_ (.A1(\channels.accum[0][5] ),
    .A2(_01360_),
    .ZN(_01382_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08915_ (.A1(_01322_),
    .A2(_01381_),
    .B(_01382_),
    .ZN(_00060_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08916_ (.I(\channels.accum[0][6] ),
    .ZN(_01383_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08917_ (.A1(_01377_),
    .A2(_01378_),
    .ZN(_01384_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _08918_ (.I(_01384_),
    .ZN(_01385_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _08919_ (.A1(_01373_),
    .A2(_01371_),
    .B(_01379_),
    .ZN(_01386_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08920_ (.A1(\channels.freq3[6] ),
    .A2(_01076_),
    .ZN(_01387_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08921_ (.A1(\channels.freq2[6] ),
    .A2(_01276_),
    .B1(_01289_),
    .B2(\channels.freq1[6] ),
    .ZN(_01388_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08922_ (.A1(_01387_),
    .A2(_01388_),
    .ZN(_01389_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _08923_ (.I0(\channels.accum[0][6] ),
    .I1(\channels.accum[1][6] ),
    .I2(\channels.accum[2][6] ),
    .I3(\channels.accum[3][6] ),
    .S0(_01147_),
    .S1(_01162_),
    .Z(_01390_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08924_ (.A1(_01389_),
    .A2(_01390_),
    .ZN(_01391_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08925_ (.I(_01391_),
    .ZN(_01392_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _08926_ (.A1(_01385_),
    .A2(_01386_),
    .A3(_01392_),
    .Z(_01393_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _08927_ (.A1(_01385_),
    .A2(_01386_),
    .B(_01392_),
    .ZN(_01394_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _08928_ (.A1(_01337_),
    .A2(_01393_),
    .A3(_01394_),
    .ZN(_01395_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08929_ (.A1(_01383_),
    .A2(_01262_),
    .B1(_01395_),
    .B2(_01318_),
    .ZN(_00061_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08930_ (.A1(_01389_),
    .A2(_01390_),
    .ZN(_01396_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08931_ (.I(_01076_),
    .Z(_01397_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08932_ (.A1(\channels.freq3[7] ),
    .A2(_01397_),
    .ZN(_01398_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08933_ (.A1(\channels.freq2[7] ),
    .A2(_01277_),
    .B1(_01289_),
    .B2(\channels.freq1[7] ),
    .ZN(_01399_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08934_ (.A1(_01398_),
    .A2(_01399_),
    .ZN(_01400_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _08935_ (.I0(\channels.accum[0][7] ),
    .I1(\channels.accum[1][7] ),
    .I2(\channels.accum[2][7] ),
    .I3(\channels.accum[3][7] ),
    .S0(_01148_),
    .S1(_01163_),
    .Z(_01401_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08936_ (.A1(_01400_),
    .A2(_01401_),
    .ZN(_01402_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _08937_ (.A1(_01396_),
    .A2(_01394_),
    .A3(_01402_),
    .Z(_01403_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _08938_ (.A1(_01396_),
    .A2(_01394_),
    .B(_01402_),
    .ZN(_01404_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08939_ (.A1(_01403_),
    .A2(_01404_),
    .ZN(_01405_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08940_ (.A1(_01349_),
    .A2(_01405_),
    .ZN(_01406_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08941_ (.A1(\channels.accum[0][7] ),
    .A2(_01360_),
    .ZN(_01407_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08942_ (.A1(_01322_),
    .A2(_01406_),
    .B(_01407_),
    .ZN(_00062_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08943_ (.I(\channels.accum[0][8] ),
    .ZN(_01408_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08944_ (.I(_01257_),
    .Z(_01409_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08945_ (.A1(_01400_),
    .A2(_01401_),
    .ZN(_01410_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _08946_ (.I(_01410_),
    .ZN(_01411_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08947_ (.A1(\channels.freq3[8] ),
    .A2(_01397_),
    .ZN(_01412_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _08948_ (.A1(\channels.freq2[8] ),
    .A2(_01277_),
    .B1(_01289_),
    .B2(\channels.freq1[8] ),
    .ZN(_01413_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08949_ (.A1(_01412_),
    .A2(_01413_),
    .ZN(_01414_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _08950_ (.I0(\channels.accum[0][8] ),
    .I1(\channels.accum[1][8] ),
    .I2(\channels.accum[2][8] ),
    .I3(\channels.accum[3][8] ),
    .S0(_01148_),
    .S1(_01163_),
    .Z(_01415_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08951_ (.A1(_01414_),
    .A2(_01415_),
    .ZN(_01416_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _08952_ (.I(_01416_),
    .ZN(_01417_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _08953_ (.A1(_01411_),
    .A2(_01404_),
    .A3(_01417_),
    .Z(_01418_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _08954_ (.A1(_01411_),
    .A2(_01404_),
    .B(_01417_),
    .ZN(_01419_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _08955_ (.A1(_01337_),
    .A2(_01418_),
    .A3(_01419_),
    .ZN(_01420_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08956_ (.I(_01254_),
    .Z(_01421_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08957_ (.A1(_01408_),
    .A2(_01409_),
    .B1(_01420_),
    .B2(_01421_),
    .ZN(_00063_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08958_ (.I(_01321_),
    .Z(_01422_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08959_ (.A1(_01414_),
    .A2(_01415_),
    .ZN(_01423_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08960_ (.A1(\channels.freq3[9] ),
    .A2(_01077_),
    .ZN(_01424_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08961_ (.I(_01276_),
    .Z(_01425_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _08962_ (.A1(\channels.freq2[9] ),
    .A2(_01425_),
    .B1(_01290_),
    .B2(\channels.freq1[9] ),
    .ZN(_01426_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08963_ (.A1(_01424_),
    .A2(_01426_),
    .ZN(_01427_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _08964_ (.I0(\channels.accum[0][9] ),
    .I1(\channels.accum[1][9] ),
    .I2(\channels.accum[2][9] ),
    .I3(\channels.accum[3][9] ),
    .S0(_01148_),
    .S1(_01163_),
    .Z(_01428_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08965_ (.A1(_01427_),
    .A2(_01428_),
    .ZN(_01429_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _08966_ (.A1(_01423_),
    .A2(_01419_),
    .A3(_01429_),
    .Z(_01430_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _08967_ (.A1(_01423_),
    .A2(_01419_),
    .B(_01429_),
    .ZN(_01431_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08968_ (.A1(_01430_),
    .A2(_01431_),
    .ZN(_01432_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08969_ (.A1(_01349_),
    .A2(_01432_),
    .ZN(_01433_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08970_ (.A1(\channels.accum[0][9] ),
    .A2(_01360_),
    .ZN(_01434_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08971_ (.A1(_01422_),
    .A2(_01433_),
    .B(_01434_),
    .ZN(_00064_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08972_ (.I(\channels.accum[0][10] ),
    .ZN(_01435_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08973_ (.I(_01298_),
    .Z(_01436_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08974_ (.A1(_01427_),
    .A2(_01428_),
    .ZN(_01437_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08975_ (.I(_01437_),
    .ZN(_01438_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08976_ (.I(_01397_),
    .Z(_01439_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08977_ (.A1(\channels.freq3[10] ),
    .A2(_01439_),
    .ZN(_01440_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _08978_ (.A1(\channels.freq2[10] ),
    .A2(_01278_),
    .B1(_01290_),
    .B2(\channels.freq1[10] ),
    .ZN(_01441_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08979_ (.A1(_01440_),
    .A2(_01441_),
    .ZN(_01442_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _08980_ (.I0(\channels.accum[0][10] ),
    .I1(\channels.accum[1][10] ),
    .I2(\channels.accum[2][10] ),
    .I3(\channels.accum[3][10] ),
    .S0(_01149_),
    .S1(_01164_),
    .Z(_01443_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08981_ (.A1(_01442_),
    .A2(_01443_),
    .ZN(_01444_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08982_ (.I(_01444_),
    .ZN(_01445_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _08983_ (.A1(_01438_),
    .A2(_01431_),
    .A3(_01445_),
    .Z(_01446_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _08984_ (.A1(_01438_),
    .A2(_01431_),
    .B(_01445_),
    .ZN(_01447_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _08985_ (.A1(_01436_),
    .A2(_01446_),
    .A3(_01447_),
    .ZN(_01448_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08986_ (.A1(_01435_),
    .A2(_01409_),
    .B1(_01448_),
    .B2(_01421_),
    .ZN(_00065_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08987_ (.I(_01299_),
    .Z(_01449_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08988_ (.A1(_01442_),
    .A2(_01443_),
    .ZN(_01450_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08989_ (.A1(\channels.freq3[11] ),
    .A2(_01079_),
    .ZN(_01451_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08990_ (.A1(\channels.freq2[11] ),
    .A2(_01279_),
    .B1(_01292_),
    .B2(\channels.freq1[11] ),
    .ZN(_01452_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08991_ (.A1(_01451_),
    .A2(_01452_),
    .ZN(_01453_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _08992_ (.I0(\channels.accum[0][11] ),
    .I1(\channels.accum[1][11] ),
    .I2(\channels.accum[2][11] ),
    .I3(\channels.accum[3][11] ),
    .S0(_01149_),
    .S1(_01165_),
    .Z(_01454_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08993_ (.A1(_01453_),
    .A2(_01454_),
    .ZN(_01455_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _08994_ (.A1(_01450_),
    .A2(_01447_),
    .A3(_01455_),
    .Z(_01456_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _08995_ (.A1(_01450_),
    .A2(_01447_),
    .B(_01455_),
    .ZN(_01457_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08996_ (.A1(_01456_),
    .A2(_01457_),
    .ZN(_01458_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08997_ (.A1(_01449_),
    .A2(_01458_),
    .ZN(_01459_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08998_ (.I(_01256_),
    .Z(_01460_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08999_ (.I(_01460_),
    .Z(_01461_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09000_ (.A1(\channels.accum[0][11] ),
    .A2(_01461_),
    .ZN(_01462_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09001_ (.A1(_01422_),
    .A2(_01459_),
    .B(_01462_),
    .ZN(_00066_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09002_ (.I(\channels.accum[0][12] ),
    .ZN(_01463_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09003_ (.A1(_01453_),
    .A2(_01454_),
    .ZN(_01464_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09004_ (.I(_01464_),
    .ZN(_01465_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09005_ (.A1(\channels.freq3[12] ),
    .A2(_01079_),
    .ZN(_01466_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09006_ (.A1(\channels.freq2[12] ),
    .A2(_01279_),
    .B1(_01292_),
    .B2(\channels.freq1[12] ),
    .ZN(_01467_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09007_ (.A1(_01466_),
    .A2(_01467_),
    .ZN(_01468_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _09008_ (.I0(\channels.accum[0][12] ),
    .I1(\channels.accum[1][12] ),
    .I2(\channels.accum[2][12] ),
    .I3(\channels.accum[3][12] ),
    .S0(_01140_),
    .S1(_01154_),
    .Z(_01469_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09009_ (.I(_01469_),
    .Z(_01470_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09010_ (.A1(_01468_),
    .A2(_01470_),
    .ZN(_01471_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09011_ (.I(_01471_),
    .ZN(_01472_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _09012_ (.A1(_01465_),
    .A2(_01457_),
    .A3(_01472_),
    .Z(_01473_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09013_ (.A1(_01465_),
    .A2(_01457_),
    .B(_01472_),
    .ZN(_01474_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _09014_ (.A1(_01436_),
    .A2(_01473_),
    .A3(_01474_),
    .ZN(_01475_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09015_ (.A1(_01463_),
    .A2(_01409_),
    .B1(_01475_),
    .B2(_01421_),
    .ZN(_00067_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09016_ (.A1(_01468_),
    .A2(_01470_),
    .ZN(_01476_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09017_ (.A1(\channels.freq3[13] ),
    .A2(_01079_),
    .ZN(_01477_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _09018_ (.A1(\channels.freq2[13] ),
    .A2(_01279_),
    .B1(_01293_),
    .B2(\channels.freq1[13] ),
    .ZN(_01478_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09019_ (.A1(_01477_),
    .A2(_01478_),
    .ZN(_01479_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09020_ (.I(_00010_),
    .Z(_01480_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _09021_ (.I0(\channels.accum[0][13] ),
    .I1(\channels.accum[1][13] ),
    .I2(\channels.accum[2][13] ),
    .I3(\channels.accum[3][13] ),
    .S0(_01138_),
    .S1(_01480_),
    .Z(_01481_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09022_ (.I(_01481_),
    .Z(_01482_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09023_ (.A1(_01479_),
    .A2(_01482_),
    .ZN(_01483_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _09024_ (.A1(_01476_),
    .A2(_01474_),
    .A3(_01483_),
    .Z(_01484_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09025_ (.A1(_01476_),
    .A2(_01474_),
    .B(_01483_),
    .ZN(_01485_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09026_ (.A1(_01484_),
    .A2(_01485_),
    .ZN(_01486_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09027_ (.A1(_01449_),
    .A2(_01486_),
    .ZN(_01487_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09028_ (.A1(\channels.accum[0][13] ),
    .A2(_01461_),
    .ZN(_01488_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09029_ (.A1(_01422_),
    .A2(_01487_),
    .B(_01488_),
    .ZN(_00068_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09030_ (.I(\channels.accum[0][14] ),
    .ZN(_01489_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09031_ (.A1(_01479_),
    .A2(_01482_),
    .ZN(_01490_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09032_ (.I(_01490_),
    .ZN(_01491_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09033_ (.A1(\channels.freq3[14] ),
    .A2(_01080_),
    .ZN(_01492_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _09034_ (.A1(\channels.freq2[14] ),
    .A2(_01280_),
    .B1(_01293_),
    .B2(\channels.freq1[14] ),
    .ZN(_01493_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09035_ (.A1(_01492_),
    .A2(_01493_),
    .ZN(_01494_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09036_ (.I(_01138_),
    .Z(_01495_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09037_ (.I(_01153_),
    .Z(_01496_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _09038_ (.I0(\channels.accum[0][14] ),
    .I1(\channels.accum[1][14] ),
    .I2(\channels.accum[2][14] ),
    .I3(\channels.accum[3][14] ),
    .S0(_01495_),
    .S1(_01496_),
    .Z(_01497_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09039_ (.I(_01497_),
    .ZN(_01498_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09040_ (.A1(_01494_),
    .A2(_01498_),
    .Z(_01499_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09041_ (.I(_01499_),
    .ZN(_01500_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _09042_ (.A1(_01491_),
    .A2(_01485_),
    .A3(_01500_),
    .Z(_01501_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09043_ (.A1(_01491_),
    .A2(_01485_),
    .B(_01500_),
    .ZN(_01502_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _09044_ (.A1(_01436_),
    .A2(_01501_),
    .A3(_01502_),
    .ZN(_01503_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09045_ (.A1(_01489_),
    .A2(_01409_),
    .B1(_01503_),
    .B2(_01421_),
    .ZN(_00069_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09046_ (.A1(_01494_),
    .A2(_01497_),
    .ZN(_01504_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09047_ (.A1(\channels.freq3[15] ),
    .A2(_01080_),
    .ZN(_01505_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _09048_ (.A1(\channels.freq2[15] ),
    .A2(_01280_),
    .B1(_01293_),
    .B2(\channels.freq1[15] ),
    .ZN(_01506_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09049_ (.A1(_01505_),
    .A2(_01506_),
    .ZN(_01507_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _09050_ (.I0(\channels.accum[0][15] ),
    .I1(\channels.accum[1][15] ),
    .I2(\channels.accum[2][15] ),
    .I3(\channels.accum[3][15] ),
    .S0(_00009_),
    .S1(_01153_),
    .Z(_01508_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09051_ (.I(_01508_),
    .ZN(_01509_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09052_ (.I(_01509_),
    .Z(_01510_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09053_ (.A1(_01507_),
    .A2(_01510_),
    .Z(_01511_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _09054_ (.A1(_01504_),
    .A2(_01502_),
    .A3(_01511_),
    .Z(_01512_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09055_ (.A1(_01504_),
    .A2(_01502_),
    .B(_01511_),
    .ZN(_01513_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09056_ (.A1(_01512_),
    .A2(_01513_),
    .ZN(_01514_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09057_ (.A1(_01449_),
    .A2(_01514_),
    .ZN(_01515_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09058_ (.A1(\channels.accum[0][15] ),
    .A2(_01461_),
    .ZN(_01516_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09059_ (.A1(_01422_),
    .A2(_01515_),
    .B(_01516_),
    .ZN(_00070_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09060_ (.I(\channels.accum[0][16] ),
    .ZN(_01517_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09061_ (.I(_01257_),
    .Z(_01518_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09062_ (.A1(_01505_),
    .A2(_01506_),
    .B(_01510_),
    .ZN(_01519_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _09063_ (.I0(\channels.accum[0][16] ),
    .I1(\channels.accum[1][16] ),
    .I2(\channels.accum[2][16] ),
    .I3(\channels.accum[3][16] ),
    .S0(_01139_),
    .S1(_01480_),
    .Z(_01520_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09064_ (.I(_01520_),
    .Z(_01521_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _09065_ (.A1(_01519_),
    .A2(_01513_),
    .A3(_01521_),
    .Z(_01522_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09066_ (.A1(_01519_),
    .A2(_01513_),
    .B(_01521_),
    .ZN(_01523_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _09067_ (.A1(_01436_),
    .A2(_01522_),
    .A3(_01523_),
    .ZN(_01524_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09068_ (.I(_01254_),
    .Z(_01525_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09069_ (.A1(_01517_),
    .A2(_01518_),
    .B1(_01524_),
    .B2(_01525_),
    .ZN(_00071_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _09070_ (.I(_01523_),
    .ZN(_01526_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _09071_ (.I0(\channels.accum[0][17] ),
    .I1(\channels.accum[1][17] ),
    .I2(\channels.accum[2][17] ),
    .I3(\channels.accum[3][17] ),
    .S0(_01139_),
    .S1(_01480_),
    .Z(_01527_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09072_ (.I(_01527_),
    .Z(_01528_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09073_ (.A1(_01526_),
    .A2(_01528_),
    .Z(_01529_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09074_ (.A1(_01323_),
    .A2(_01529_),
    .Z(_01530_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09075_ (.A1(\channels.accum[0][17] ),
    .A2(_01334_),
    .B1(_01530_),
    .B2(_01255_),
    .ZN(_01531_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09076_ (.I(_01531_),
    .ZN(_00072_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09077_ (.I(\channels.accum[0][18] ),
    .ZN(_01532_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _09078_ (.I0(\channels.accum[0][18] ),
    .I1(\channels.accum[1][18] ),
    .I2(\channels.accum[2][18] ),
    .I3(\channels.accum[3][18] ),
    .S0(_01495_),
    .S1(_01496_),
    .Z(_01533_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09079_ (.I(_01533_),
    .Z(_01534_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09080_ (.A1(_01526_),
    .A2(_01528_),
    .B(_01534_),
    .ZN(_01535_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09081_ (.A1(_01526_),
    .A2(_01528_),
    .A3(_01534_),
    .ZN(_01536_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09082_ (.I(_01536_),
    .Z(_01537_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09083_ (.A1(_01323_),
    .A2(_01537_),
    .ZN(_01538_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09084_ (.A1(_01535_),
    .A2(_01538_),
    .Z(_01539_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09085_ (.A1(_01532_),
    .A2(_01518_),
    .B1(_01539_),
    .B2(_01525_),
    .ZN(_00073_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09086_ (.I(_01321_),
    .Z(_01540_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _09087_ (.I0(\channels.accum[0][19] ),
    .I1(\channels.accum[1][19] ),
    .I2(\channels.accum[2][19] ),
    .I3(\channels.accum[3][19] ),
    .S0(_01495_),
    .S1(_01496_),
    .Z(_01541_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09088_ (.I(_01541_),
    .Z(_01542_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _09089_ (.I(_01542_),
    .ZN(_01543_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09090_ (.A1(_01537_),
    .A2(_01543_),
    .Z(_01544_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09091_ (.A1(_01449_),
    .A2(_01544_),
    .ZN(_01545_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09092_ (.A1(\channels.accum[0][19] ),
    .A2(_01461_),
    .ZN(_01546_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09093_ (.A1(_01540_),
    .A2(_01545_),
    .B(_01546_),
    .ZN(_00074_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09094_ (.I(\channels.accum[0][20] ),
    .ZN(_01547_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09095_ (.A1(_01537_),
    .A2(_01543_),
    .ZN(_01548_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _09096_ (.I0(\channels.accum[0][20] ),
    .I1(\channels.accum[1][20] ),
    .I2(\channels.accum[2][20] ),
    .I3(\channels.accum[3][20] ),
    .S0(_01138_),
    .S1(_01153_),
    .Z(_01549_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09097_ (.I(_01549_),
    .Z(_01550_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09098_ (.A1(_01548_),
    .A2(_01550_),
    .Z(_01551_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09099_ (.A1(_01300_),
    .A2(_01551_),
    .ZN(_01552_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09100_ (.A1(_01547_),
    .A2(_01518_),
    .B1(_01552_),
    .B2(_01525_),
    .ZN(_00075_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _09101_ (.I(_01549_),
    .ZN(_01553_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _09102_ (.A1(_01536_),
    .A2(_01543_),
    .A3(_01553_),
    .ZN(_01554_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _09103_ (.I0(\channels.accum[0][21] ),
    .I1(\channels.accum[1][21] ),
    .I2(\channels.accum[2][21] ),
    .I3(\channels.accum[3][21] ),
    .S0(_01139_),
    .S1(_01480_),
    .Z(_01555_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09104_ (.I(_01555_),
    .Z(_01556_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09105_ (.A1(_01554_),
    .A2(_01556_),
    .Z(_01557_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09106_ (.A1(_01554_),
    .A2(_01556_),
    .ZN(_01558_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _09107_ (.A1(_01323_),
    .A2(_01557_),
    .A3(_01558_),
    .ZN(_01559_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09108_ (.I(_01460_),
    .Z(_01560_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09109_ (.A1(\channels.accum[0][21] ),
    .A2(_01560_),
    .ZN(_01561_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09110_ (.A1(_01540_),
    .A2(_01559_),
    .B(_01561_),
    .ZN(_00076_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09111_ (.I(\channels.accum[0][22] ),
    .ZN(_01562_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09112_ (.I(\channels.accum[1][22] ),
    .ZN(_01563_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09113_ (.I(\channels.accum[2][22] ),
    .ZN(_01564_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09114_ (.I(\channels.accum[3][22] ),
    .ZN(_01565_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _09115_ (.I0(_01562_),
    .I1(_01563_),
    .I2(_01564_),
    .I3(_01565_),
    .S0(_01140_),
    .S1(_01154_),
    .Z(_01566_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09116_ (.A1(_01558_),
    .A2(_01566_),
    .Z(_01567_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09117_ (.A1(_01300_),
    .A2(_01567_),
    .ZN(_01568_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09118_ (.A1(_01562_),
    .A2(_01518_),
    .B1(_01568_),
    .B2(_01525_),
    .ZN(_00077_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09119_ (.A1(_01558_),
    .A2(_01566_),
    .ZN(_01569_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09120_ (.A1(_01086_),
    .A2(_01569_),
    .Z(_01570_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09121_ (.A1(_01300_),
    .A2(_01570_),
    .ZN(_01571_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09122_ (.A1(\channels.accum[0][23] ),
    .A2(_01560_),
    .ZN(_01572_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09123_ (.A1(_01540_),
    .A2(_01571_),
    .B(_01572_),
    .ZN(_00078_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09124_ (.I(\channels.lfsr[0][17] ),
    .ZN(_01573_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09125_ (.I(\channels.lfsr[1][17] ),
    .ZN(_01574_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09126_ (.I(\channels.lfsr[2][17] ),
    .ZN(_01575_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09127_ (.I(\channels.lfsr[3][17] ),
    .ZN(_01576_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _09128_ (.I0(_01573_),
    .I1(_01574_),
    .I2(_01575_),
    .I3(_01576_),
    .S0(_01201_),
    .S1(_01304_),
    .Z(_01577_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _09129_ (.I0(\channels.lfsr[0][22] ),
    .I1(\channels.lfsr[1][22] ),
    .I2(\channels.lfsr[2][22] ),
    .I3(\channels.lfsr[3][22] ),
    .S0(_01201_),
    .S1(_01304_),
    .Z(_01578_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09130_ (.A1(_01577_),
    .A2(_01578_),
    .ZN(_01579_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09131_ (.A1(_01270_),
    .A2(_01579_),
    .ZN(_01580_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09132_ (.I(_01082_),
    .Z(_01581_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09133_ (.I(_01249_),
    .Z(_01582_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _09134_ (.I(_01582_),
    .Z(_01583_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _09135_ (.A1(_01583_),
    .A2(_01264_),
    .B(_01095_),
    .ZN(_01584_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09136_ (.I(_01584_),
    .Z(_01585_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09137_ (.I(_01585_),
    .ZN(_01586_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _09138_ (.A1(_01270_),
    .A2(_01537_),
    .A3(_01542_),
    .A4(_01586_),
    .ZN(_01587_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _09139_ (.A1(_01581_),
    .A2(_01587_),
    .Z(_01588_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09140_ (.I(_01588_),
    .Z(_01589_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09141_ (.A1(_01043_),
    .A2(_01588_),
    .ZN(_01590_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09142_ (.I(_01590_),
    .Z(_01591_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09143_ (.I(_01591_),
    .Z(_01592_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09144_ (.I(\channels.lfsr[2][0] ),
    .ZN(_01593_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09145_ (.A1(_01580_),
    .A2(_01589_),
    .B1(_01592_),
    .B2(_01593_),
    .ZN(_00079_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09146_ (.I(\channels.lfsr[2][1] ),
    .ZN(_01594_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09147_ (.I(\channels.lfsr[0][0] ),
    .ZN(_01595_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09148_ (.I(\channels.lfsr[1][0] ),
    .ZN(_01596_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09149_ (.I(\channels.lfsr[3][0] ),
    .ZN(_01597_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _09150_ (.I0(_01595_),
    .I1(_01596_),
    .I2(_01593_),
    .I3(_01597_),
    .S0(_01140_),
    .S1(_01154_),
    .Z(_01598_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09151_ (.I(_01589_),
    .Z(_01599_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09152_ (.A1(_01594_),
    .A2(_01592_),
    .B1(_01598_),
    .B2(_01599_),
    .ZN(_00080_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09153_ (.I(\channels.lfsr[2][2] ),
    .ZN(_01600_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09154_ (.I(\channels.lfsr[0][1] ),
    .ZN(_01601_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09155_ (.I(\channels.lfsr[1][1] ),
    .ZN(_01602_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09156_ (.I(\channels.lfsr[3][1] ),
    .ZN(_01603_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09157_ (.I(_01201_),
    .Z(_01604_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09158_ (.I(_01604_),
    .Z(_01605_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09159_ (.I(_01304_),
    .Z(_01606_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09160_ (.I(_01606_),
    .Z(_01607_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _09161_ (.I0(_01601_),
    .I1(_01602_),
    .I2(_01594_),
    .I3(_01603_),
    .S0(_01605_),
    .S1(_01607_),
    .Z(_01608_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09162_ (.A1(_01600_),
    .A2(_01592_),
    .B1(_01608_),
    .B2(_01599_),
    .ZN(_00081_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09163_ (.I(\channels.lfsr[2][3] ),
    .ZN(_01609_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09164_ (.I(_01590_),
    .Z(_01610_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09165_ (.I(_01610_),
    .Z(_01611_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09166_ (.I(\channels.lfsr[0][2] ),
    .ZN(_01612_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09167_ (.I(\channels.lfsr[1][2] ),
    .ZN(_01613_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09168_ (.I(\channels.lfsr[3][2] ),
    .ZN(_01614_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _09169_ (.I0(_01612_),
    .I1(_01613_),
    .I2(_01600_),
    .I3(_01614_),
    .S0(_01141_),
    .S1(_01155_),
    .Z(_01615_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09170_ (.A1(_01609_),
    .A2(_01611_),
    .B1(_01615_),
    .B2(_01599_),
    .ZN(_00082_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09171_ (.I(\channels.lfsr[2][4] ),
    .ZN(_01616_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09172_ (.I(\channels.lfsr[0][3] ),
    .ZN(_01617_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09173_ (.I(\channels.lfsr[1][3] ),
    .ZN(_01618_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09174_ (.I(\channels.lfsr[3][3] ),
    .ZN(_01619_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _09175_ (.I0(_01617_),
    .I1(_01618_),
    .I2(_01609_),
    .I3(_01619_),
    .S0(_01605_),
    .S1(_01607_),
    .Z(_01620_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09176_ (.A1(_01616_),
    .A2(_01611_),
    .B1(_01620_),
    .B2(_01599_),
    .ZN(_00083_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09177_ (.I(\channels.lfsr[2][5] ),
    .ZN(_01621_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09178_ (.I(\channels.lfsr[0][4] ),
    .ZN(_01622_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09179_ (.I(\channels.lfsr[1][4] ),
    .ZN(_01623_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09180_ (.I(\channels.lfsr[3][4] ),
    .ZN(_01624_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _09181_ (.I0(_01622_),
    .I1(_01623_),
    .I2(_01616_),
    .I3(_01624_),
    .S0(_01605_),
    .S1(_01607_),
    .Z(_01625_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09182_ (.I(_01588_),
    .Z(_01626_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09183_ (.I(_01626_),
    .Z(_01627_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09184_ (.A1(_01621_),
    .A2(_01611_),
    .B1(_01625_),
    .B2(_01627_),
    .ZN(_00084_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09185_ (.I(\channels.lfsr[2][6] ),
    .ZN(_01628_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09186_ (.I(\channels.lfsr[0][5] ),
    .ZN(_01629_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09187_ (.I(\channels.lfsr[1][5] ),
    .ZN(_01630_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09188_ (.I(\channels.lfsr[3][5] ),
    .ZN(_01631_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _09189_ (.I0(_01629_),
    .I1(_01630_),
    .I2(_01621_),
    .I3(_01631_),
    .S0(_01141_),
    .S1(_01155_),
    .Z(_01632_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09190_ (.A1(_01628_),
    .A2(_01611_),
    .B1(_01632_),
    .B2(_01627_),
    .ZN(_00085_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09191_ (.I(\channels.lfsr[2][7] ),
    .ZN(_01633_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09192_ (.I(_01610_),
    .Z(_01634_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09193_ (.I(\channels.lfsr[0][6] ),
    .ZN(_01635_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09194_ (.I(\channels.lfsr[1][6] ),
    .ZN(_01636_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09195_ (.I(\channels.lfsr[3][6] ),
    .ZN(_01637_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _09196_ (.I0(_01635_),
    .I1(_01636_),
    .I2(_01628_),
    .I3(_01637_),
    .S0(_01605_),
    .S1(_01607_),
    .Z(_01638_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09197_ (.A1(_01633_),
    .A2(_01634_),
    .B1(_01638_),
    .B2(_01627_),
    .ZN(_00086_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09198_ (.I(\channels.lfsr[2][8] ),
    .ZN(_01639_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09199_ (.I(\channels.lfsr[0][7] ),
    .ZN(_01640_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09200_ (.I(\channels.lfsr[1][7] ),
    .ZN(_01641_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09201_ (.I(\channels.lfsr[3][7] ),
    .ZN(_01642_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09202_ (.I(_01604_),
    .Z(_01643_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09203_ (.I(_01606_),
    .Z(_01644_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _09204_ (.I0(_01640_),
    .I1(_01641_),
    .I2(_01633_),
    .I3(_01642_),
    .S0(_01643_),
    .S1(_01644_),
    .Z(_01645_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09205_ (.A1(_01639_),
    .A2(_01634_),
    .B1(_01645_),
    .B2(_01627_),
    .ZN(_00087_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09206_ (.I(\channels.lfsr[2][9] ),
    .ZN(_01646_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09207_ (.I(\channels.lfsr[0][8] ),
    .ZN(_01647_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09208_ (.I(\channels.lfsr[1][8] ),
    .ZN(_01648_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09209_ (.I(\channels.lfsr[3][8] ),
    .ZN(_01649_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _09210_ (.I0(_01647_),
    .I1(_01648_),
    .I2(_01639_),
    .I3(_01649_),
    .S0(_01643_),
    .S1(_01644_),
    .Z(_01650_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09211_ (.I(_01626_),
    .Z(_01651_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09212_ (.A1(_01646_),
    .A2(_01634_),
    .B1(_01650_),
    .B2(_01651_),
    .ZN(_00088_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09213_ (.I(\channels.lfsr[2][10] ),
    .ZN(_01652_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09214_ (.I(\channels.lfsr[0][9] ),
    .ZN(_01653_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09215_ (.I(\channels.lfsr[1][9] ),
    .ZN(_01654_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09216_ (.I(\channels.lfsr[3][9] ),
    .ZN(_01655_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09217_ (.I(_01155_),
    .Z(_01656_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _09218_ (.I0(_01653_),
    .I1(_01654_),
    .I2(_01646_),
    .I3(_01655_),
    .S0(_01142_),
    .S1(_01656_),
    .Z(_01657_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09219_ (.A1(_01652_),
    .A2(_01634_),
    .B1(_01657_),
    .B2(_01651_),
    .ZN(_00089_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09220_ (.I(\channels.lfsr[2][11] ),
    .ZN(_01658_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09221_ (.I(_01610_),
    .Z(_01659_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09222_ (.I(\channels.lfsr[0][10] ),
    .ZN(_01660_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09223_ (.I(\channels.lfsr[1][10] ),
    .ZN(_01661_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09224_ (.I(\channels.lfsr[3][10] ),
    .ZN(_01662_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _09225_ (.I0(_01660_),
    .I1(_01661_),
    .I2(_01652_),
    .I3(_01662_),
    .S0(_01643_),
    .S1(_01644_),
    .Z(_01663_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09226_ (.A1(_01658_),
    .A2(_01659_),
    .B1(_01663_),
    .B2(_01651_),
    .ZN(_00090_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09227_ (.I(\channels.lfsr[2][12] ),
    .ZN(_01664_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09228_ (.I(\channels.lfsr[0][11] ),
    .ZN(_01665_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09229_ (.I(\channels.lfsr[1][11] ),
    .ZN(_01666_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09230_ (.I(\channels.lfsr[3][11] ),
    .ZN(_01667_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _09231_ (.I0(_01665_),
    .I1(_01666_),
    .I2(_01658_),
    .I3(_01667_),
    .S0(_01305_),
    .S1(_01656_),
    .Z(_01668_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09232_ (.A1(_01664_),
    .A2(_01659_),
    .B1(_01668_),
    .B2(_01651_),
    .ZN(_00091_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09233_ (.I(\channels.lfsr[2][13] ),
    .ZN(_01669_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09234_ (.I(\channels.lfsr[0][12] ),
    .ZN(_01670_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09235_ (.I(\channels.lfsr[1][12] ),
    .ZN(_01671_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09236_ (.I(\channels.lfsr[3][12] ),
    .ZN(_01672_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _09237_ (.I0(_01670_),
    .I1(_01671_),
    .I2(_01664_),
    .I3(_01672_),
    .S0(_01643_),
    .S1(_01644_),
    .Z(_01673_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09238_ (.I(_01626_),
    .Z(_01674_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09239_ (.A1(_01669_),
    .A2(_01659_),
    .B1(_01673_),
    .B2(_01674_),
    .ZN(_00092_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09240_ (.I(\channels.lfsr[2][14] ),
    .ZN(_01675_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09241_ (.I(\channels.lfsr[0][13] ),
    .ZN(_01676_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09242_ (.I(\channels.lfsr[1][13] ),
    .ZN(_01677_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09243_ (.I(\channels.lfsr[3][13] ),
    .ZN(_01678_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09244_ (.I(_01604_),
    .Z(_01679_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09245_ (.I(_01606_),
    .Z(_01680_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _09246_ (.I0(_01676_),
    .I1(_01677_),
    .I2(_01669_),
    .I3(_01678_),
    .S0(_01679_),
    .S1(_01680_),
    .Z(_01681_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09247_ (.A1(_01675_),
    .A2(_01659_),
    .B1(_01681_),
    .B2(_01674_),
    .ZN(_00093_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09248_ (.I(\channels.lfsr[2][15] ),
    .ZN(_01682_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09249_ (.I(_01610_),
    .Z(_01683_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09250_ (.I(\channels.lfsr[0][14] ),
    .ZN(_01684_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09251_ (.I(\channels.lfsr[1][14] ),
    .ZN(_01685_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09252_ (.I(\channels.lfsr[3][14] ),
    .ZN(_01686_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09253_ (.I(_01656_),
    .Z(_01687_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09254_ (.I(_01687_),
    .Z(_01688_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _09255_ (.I0(_01684_),
    .I1(_01685_),
    .I2(_01675_),
    .I3(_01686_),
    .S0(_01144_),
    .S1(_01688_),
    .Z(_01689_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09256_ (.A1(_01682_),
    .A2(_01683_),
    .B1(_01689_),
    .B2(_01674_),
    .ZN(_00094_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09257_ (.I(\channels.lfsr[2][16] ),
    .ZN(_01690_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09258_ (.I(\channels.lfsr[0][15] ),
    .ZN(_01691_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09259_ (.I(\channels.lfsr[1][15] ),
    .ZN(_01692_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09260_ (.I(\channels.lfsr[3][15] ),
    .ZN(_01693_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _09261_ (.I0(_01691_),
    .I1(_01692_),
    .I2(_01682_),
    .I3(_01693_),
    .S0(_01679_),
    .S1(_01680_),
    .Z(_01694_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09262_ (.A1(_01690_),
    .A2(_01683_),
    .B1(_01694_),
    .B2(_01674_),
    .ZN(_00095_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09263_ (.I(\channels.lfsr[0][16] ),
    .ZN(_01695_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09264_ (.I(\channels.lfsr[1][16] ),
    .ZN(_01696_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09265_ (.I(\channels.lfsr[3][16] ),
    .ZN(_01697_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _09266_ (.I0(_01695_),
    .I1(_01696_),
    .I2(_01690_),
    .I3(_01697_),
    .S0(_01679_),
    .S1(_01680_),
    .Z(_01698_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09267_ (.I(_01626_),
    .Z(_01699_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09268_ (.A1(_01575_),
    .A2(_01683_),
    .B1(_01698_),
    .B2(_01699_),
    .ZN(_00096_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09269_ (.I(\channels.lfsr[2][18] ),
    .ZN(_01700_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09270_ (.A1(_01577_),
    .A2(_01589_),
    .B1(_01592_),
    .B2(_01700_),
    .ZN(_00097_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09271_ (.I(\channels.lfsr[2][19] ),
    .ZN(_01701_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09272_ (.I(\channels.lfsr[0][18] ),
    .ZN(_01702_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09273_ (.I(\channels.lfsr[1][18] ),
    .ZN(_01703_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09274_ (.I(\channels.lfsr[3][18] ),
    .ZN(_01704_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _09275_ (.I0(_01702_),
    .I1(_01703_),
    .I2(_01700_),
    .I3(_01704_),
    .S0(_01144_),
    .S1(_01158_),
    .Z(_01705_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09276_ (.A1(_01701_),
    .A2(_01683_),
    .B1(_01705_),
    .B2(_01699_),
    .ZN(_00098_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09277_ (.I(\channels.lfsr[2][20] ),
    .ZN(_01706_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09278_ (.I(\channels.lfsr[0][19] ),
    .ZN(_01707_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09279_ (.I(\channels.lfsr[1][19] ),
    .ZN(_01708_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09280_ (.I(\channels.lfsr[3][19] ),
    .ZN(_01709_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _09281_ (.I0(_01707_),
    .I1(_01708_),
    .I2(_01701_),
    .I3(_01709_),
    .S0(_01679_),
    .S1(_01680_),
    .Z(_01710_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09282_ (.A1(_01706_),
    .A2(_01591_),
    .B1(_01710_),
    .B2(_01699_),
    .ZN(_00099_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09283_ (.I(\channels.lfsr[2][21] ),
    .ZN(_01711_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09284_ (.I(\channels.lfsr[0][20] ),
    .ZN(_01712_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09285_ (.I(\channels.lfsr[1][20] ),
    .ZN(_01713_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09286_ (.I(\channels.lfsr[3][20] ),
    .ZN(_01714_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _09287_ (.I0(_01712_),
    .I1(_01713_),
    .I2(_01706_),
    .I3(_01714_),
    .S0(_01145_),
    .S1(_01328_),
    .Z(_01715_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09288_ (.A1(_01711_),
    .A2(_01591_),
    .B1(_01715_),
    .B2(_01699_),
    .ZN(_00100_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09289_ (.I(\channels.lfsr[2][22] ),
    .ZN(_01716_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09290_ (.I(\channels.lfsr[0][21] ),
    .ZN(_01717_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09291_ (.I(\channels.lfsr[1][21] ),
    .ZN(_01718_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09292_ (.I(\channels.lfsr[3][21] ),
    .ZN(_01719_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _09293_ (.I0(_01717_),
    .I1(_01718_),
    .I2(_01711_),
    .I3(_01719_),
    .S0(_01604_),
    .S1(_01606_),
    .Z(_01720_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09294_ (.A1(_01716_),
    .A2(_01591_),
    .B1(_01720_),
    .B2(_01589_),
    .ZN(_00101_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _09295_ (.A1(_01282_),
    .A2(_01587_),
    .Z(_01721_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09296_ (.I(_01721_),
    .Z(_01722_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09297_ (.I(_01722_),
    .Z(_01723_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _09298_ (.I(_01032_),
    .Z(_01724_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09299_ (.A1(_01724_),
    .A2(_01721_),
    .ZN(_01725_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09300_ (.I(_01725_),
    .Z(_01726_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09301_ (.I(_01726_),
    .Z(_01727_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09302_ (.A1(_01580_),
    .A2(_01723_),
    .B1(_01727_),
    .B2(_01596_),
    .ZN(_00102_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09303_ (.A1(_01598_),
    .A2(_01723_),
    .B1(_01727_),
    .B2(_01602_),
    .ZN(_00103_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09304_ (.A1(_01608_),
    .A2(_01723_),
    .B1(_01727_),
    .B2(_01613_),
    .ZN(_00104_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09305_ (.A1(_01615_),
    .A2(_01723_),
    .B1(_01727_),
    .B2(_01618_),
    .ZN(_00105_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09306_ (.I(_01721_),
    .Z(_01728_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09307_ (.I(_01728_),
    .Z(_01729_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09308_ (.I(_01725_),
    .Z(_01730_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09309_ (.I(_01730_),
    .Z(_01731_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09310_ (.A1(_01620_),
    .A2(_01729_),
    .B1(_01731_),
    .B2(_01623_),
    .ZN(_00106_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09311_ (.A1(_01625_),
    .A2(_01729_),
    .B1(_01731_),
    .B2(_01630_),
    .ZN(_00107_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09312_ (.A1(_01632_),
    .A2(_01729_),
    .B1(_01731_),
    .B2(_01636_),
    .ZN(_00108_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09313_ (.A1(_01638_),
    .A2(_01729_),
    .B1(_01731_),
    .B2(_01641_),
    .ZN(_00109_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09314_ (.I(_01728_),
    .Z(_01732_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09315_ (.I(_01730_),
    .Z(_01733_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09316_ (.A1(_01645_),
    .A2(_01732_),
    .B1(_01733_),
    .B2(_01648_),
    .ZN(_00110_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09317_ (.A1(_01650_),
    .A2(_01732_),
    .B1(_01733_),
    .B2(_01654_),
    .ZN(_00111_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09318_ (.A1(_01657_),
    .A2(_01732_),
    .B1(_01733_),
    .B2(_01661_),
    .ZN(_00112_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09319_ (.A1(_01663_),
    .A2(_01732_),
    .B1(_01733_),
    .B2(_01666_),
    .ZN(_00113_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09320_ (.I(_01728_),
    .Z(_01734_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09321_ (.I(_01730_),
    .Z(_01735_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09322_ (.A1(_01668_),
    .A2(_01734_),
    .B1(_01735_),
    .B2(_01671_),
    .ZN(_00114_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09323_ (.A1(_01673_),
    .A2(_01734_),
    .B1(_01735_),
    .B2(_01677_),
    .ZN(_00115_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09324_ (.A1(_01681_),
    .A2(_01734_),
    .B1(_01735_),
    .B2(_01685_),
    .ZN(_00116_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09325_ (.A1(_01689_),
    .A2(_01734_),
    .B1(_01735_),
    .B2(_01692_),
    .ZN(_00117_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09326_ (.I(_01728_),
    .Z(_01736_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09327_ (.I(_01730_),
    .Z(_01737_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09328_ (.A1(_01694_),
    .A2(_01736_),
    .B1(_01737_),
    .B2(_01696_),
    .ZN(_00118_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09329_ (.A1(_01698_),
    .A2(_01736_),
    .B1(_01737_),
    .B2(_01574_),
    .ZN(_00119_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09330_ (.A1(_01577_),
    .A2(_01736_),
    .B1(_01737_),
    .B2(_01703_),
    .ZN(_00120_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09331_ (.A1(_01705_),
    .A2(_01736_),
    .B1(_01737_),
    .B2(_01708_),
    .ZN(_00121_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09332_ (.A1(_01710_),
    .A2(_01722_),
    .B1(_01726_),
    .B2(_01713_),
    .ZN(_00122_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09333_ (.A1(_01715_),
    .A2(_01722_),
    .B1(_01726_),
    .B2(_01718_),
    .ZN(_00123_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09334_ (.I(\channels.lfsr[1][22] ),
    .ZN(_01738_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09335_ (.A1(_01720_),
    .A2(_01722_),
    .B1(_01726_),
    .B2(_01738_),
    .ZN(_00124_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09336_ (.I(net8),
    .ZN(_01739_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09337_ (.I(_01739_),
    .Z(_01740_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09338_ (.I(_01740_),
    .Z(_01741_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09339_ (.I(_01741_),
    .Z(_01742_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09340_ (.I(_01013_),
    .Z(_01743_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09341_ (.I(\filters.filt_1 ),
    .Z(_01744_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09342_ (.I(_01744_),
    .Z(_01745_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09343_ (.I(_01745_),
    .Z(_01746_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09344_ (.I(_01746_),
    .Z(_01747_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _09345_ (.I(_01747_),
    .Z(_01748_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09346_ (.I(_01013_),
    .Z(_01749_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09347_ (.I(_01062_),
    .Z(_01750_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09348_ (.I(_01750_),
    .Z(_01751_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09349_ (.I(_01751_),
    .Z(_01752_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09350_ (.I(_01752_),
    .Z(_01753_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09351_ (.A1(_01748_),
    .A2(_01749_),
    .B(_01753_),
    .ZN(_01754_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09352_ (.A1(_01742_),
    .A2(_01743_),
    .B(_01754_),
    .ZN(_00125_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _09353_ (.I(net9),
    .ZN(_01755_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09354_ (.I(_01755_),
    .Z(_01756_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09355_ (.I(_01756_),
    .Z(_01757_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09356_ (.I(\filters.filt_2 ),
    .Z(_01758_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09357_ (.I(_01758_),
    .Z(_01759_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09358_ (.I(_01759_),
    .Z(_01760_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09359_ (.I(_01760_),
    .Z(_01761_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _09360_ (.I(_01761_),
    .Z(_01762_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09361_ (.I(_01752_),
    .Z(_01763_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09362_ (.A1(_01762_),
    .A2(_01749_),
    .B(_01763_),
    .ZN(_01764_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09363_ (.A1(_01757_),
    .A2(_01743_),
    .B(_01764_),
    .ZN(_00126_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _09364_ (.I(net10),
    .ZN(_01765_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09365_ (.I(_01765_),
    .Z(_01766_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09366_ (.I(_01766_),
    .Z(_01767_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09367_ (.I(\filters.filt_3 ),
    .Z(_01768_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09368_ (.I(_01768_),
    .Z(_01769_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09369_ (.I(_01769_),
    .Z(_01770_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09370_ (.I(_01770_),
    .Z(_01771_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09371_ (.I(_01771_),
    .Z(_01772_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09372_ (.I(_01772_),
    .Z(_01773_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09373_ (.A1(_01773_),
    .A2(_01749_),
    .B(_01763_),
    .ZN(_01774_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09374_ (.A1(_01767_),
    .A2(_01743_),
    .B(_01774_),
    .ZN(_00127_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09375_ (.I(net11),
    .ZN(_01775_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09376_ (.I(_01775_),
    .Z(_01776_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09377_ (.I(_01776_),
    .Z(_01777_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09378_ (.A1(\filters.res_filt[3] ),
    .A2(_01749_),
    .B(_01763_),
    .ZN(_01778_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09379_ (.A1(_01777_),
    .A2(_01743_),
    .B(_01778_),
    .ZN(_00128_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09380_ (.I(_01003_),
    .Z(_01779_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09381_ (.I(_01779_),
    .Z(_01780_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09382_ (.I(_01780_),
    .Z(_01781_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09383_ (.I(net6),
    .ZN(_01782_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09384_ (.A1(_01782_),
    .A2(net5),
    .ZN(_01783_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _09385_ (.I(net3),
    .ZN(_01784_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09386_ (.A1(net4),
    .A2(_01784_),
    .ZN(_01785_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _09387_ (.I(net2),
    .ZN(_01786_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _09388_ (.I(net1),
    .ZN(_01787_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09389_ (.A1(_01786_),
    .A2(_01787_),
    .ZN(_01788_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09390_ (.I(_01788_),
    .Z(_01789_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _09391_ (.A1(_01783_),
    .A2(_01785_),
    .A3(_01789_),
    .ZN(_01790_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09392_ (.I(_01790_),
    .Z(_01791_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09393_ (.A1(_01781_),
    .A2(_01791_),
    .Z(_01792_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09394_ (.I(_01792_),
    .Z(_01793_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09395_ (.I(_01792_),
    .Z(_01794_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09396_ (.A1(\filters.mode_vol[0] ),
    .A2(_01794_),
    .B(_01763_),
    .ZN(_01795_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09397_ (.A1(_01742_),
    .A2(_01793_),
    .B(_01795_),
    .ZN(_00133_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09398_ (.I(_01752_),
    .Z(_01796_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09399_ (.A1(\filters.mode_vol[1] ),
    .A2(_01794_),
    .B(_01796_),
    .ZN(_01797_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09400_ (.A1(_01757_),
    .A2(_01793_),
    .B(_01797_),
    .ZN(_00134_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09401_ (.A1(\filters.mode_vol[2] ),
    .A2(_01794_),
    .B(_01796_),
    .ZN(_01798_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09402_ (.A1(_01767_),
    .A2(_01793_),
    .B(_01798_),
    .ZN(_00135_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09403_ (.A1(\filters.mode_vol[3] ),
    .A2(_01794_),
    .B(_01796_),
    .ZN(_01799_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09404_ (.A1(_01777_),
    .A2(_01793_),
    .B(_01799_),
    .ZN(_00136_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09405_ (.I(_01017_),
    .Z(_01800_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09406_ (.I(_01800_),
    .Z(_01801_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09407_ (.I(_01792_),
    .Z(_01802_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09408_ (.I(_01792_),
    .Z(_01803_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09409_ (.A1(\filters.lp ),
    .A2(_01803_),
    .B(_01796_),
    .ZN(_01804_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09410_ (.A1(_01801_),
    .A2(_01802_),
    .B(_01804_),
    .ZN(_00137_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09411_ (.I(_01006_),
    .Z(_01805_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09412_ (.I(_01805_),
    .Z(_01806_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09413_ (.I(_01806_),
    .Z(_01807_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09414_ (.I(_01751_),
    .Z(_01808_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09415_ (.I(_01808_),
    .Z(_01809_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09416_ (.A1(\filters.bp ),
    .A2(_01803_),
    .B(_01809_),
    .ZN(_01810_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09417_ (.A1(_01807_),
    .A2(_01802_),
    .B(_01810_),
    .ZN(_00138_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09418_ (.I(net14),
    .Z(_01811_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _09419_ (.I(_01811_),
    .ZN(_01812_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09420_ (.I(_01812_),
    .Z(_01813_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09421_ (.I(_01813_),
    .Z(_01814_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09422_ (.A1(\filters.hp ),
    .A2(_01803_),
    .B(_01809_),
    .ZN(_01815_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09423_ (.A1(_01814_),
    .A2(_01802_),
    .B(_01815_),
    .ZN(_00139_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _09424_ (.I(net15),
    .ZN(_01816_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09425_ (.I(_01816_),
    .Z(_01817_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09426_ (.I(_01817_),
    .Z(_01818_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09427_ (.I(_01818_),
    .Z(_01819_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09428_ (.A1(\filters.mode_vol[7] ),
    .A2(_01803_),
    .B(_01809_),
    .ZN(_01820_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09429_ (.A1(_01819_),
    .A2(_01802_),
    .B(_01820_),
    .ZN(_00140_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09430_ (.I(_01102_),
    .Z(_01821_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09431_ (.I(_01821_),
    .Z(_01822_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09432_ (.I(_01822_),
    .Z(_01823_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09433_ (.I(_01001_),
    .Z(_01824_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09434_ (.I(_01824_),
    .Z(_01825_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09435_ (.I(_01785_),
    .Z(_01826_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09436_ (.A1(_01782_),
    .A2(_00998_),
    .ZN(_01827_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09437_ (.I(_01827_),
    .Z(_01828_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _09438_ (.A1(_01825_),
    .A2(_01826_),
    .A3(_01828_),
    .ZN(_01829_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09439_ (.I(_01829_),
    .Z(_01830_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09440_ (.A1(net4),
    .A2(net3),
    .ZN(_01831_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09441_ (.I(_01831_),
    .Z(_01832_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _09442_ (.A1(_01825_),
    .A2(_01828_),
    .A3(_01832_),
    .ZN(_01833_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09443_ (.I(_01833_),
    .Z(_01834_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09444_ (.A1(\channels.ctrl_reg2[0] ),
    .A2(_01830_),
    .B1(_01834_),
    .B2(\channels.freq3[8] ),
    .ZN(_01835_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09445_ (.I(_01788_),
    .Z(_01836_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _09446_ (.A1(_01836_),
    .A2(_01828_),
    .A3(_01832_),
    .ZN(_01837_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09447_ (.I(_01837_),
    .Z(_01838_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09448_ (.A1(_01786_),
    .A2(net1),
    .ZN(_01839_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _09449_ (.A1(_00997_),
    .A2(_01784_),
    .A3(_00999_),
    .ZN(_01840_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09450_ (.A1(_01839_),
    .A2(_01840_),
    .ZN(_01841_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09451_ (.I(_01841_),
    .Z(_01842_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09452_ (.A1(\channels.atk_dec2[0] ),
    .A2(_01838_),
    .B1(_01842_),
    .B2(\channels.pw3[8] ),
    .ZN(_01843_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09453_ (.I(_01002_),
    .Z(_01844_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09454_ (.A1(net6),
    .A2(net5),
    .ZN(_01845_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _09455_ (.A1(_01786_),
    .A2(net1),
    .A3(_01845_),
    .ZN(_01846_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09456_ (.A1(_01826_),
    .A2(_01846_),
    .ZN(_01847_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09457_ (.I(_01847_),
    .Z(_01848_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09458_ (.A1(_01000_),
    .A2(_01839_),
    .ZN(_01849_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09459_ (.A1(net2),
    .A2(_01787_),
    .ZN(_01850_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09460_ (.A1(_01000_),
    .A2(_01850_),
    .ZN(_01851_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _09461_ (.A1(\filters.cutoff_lut[6] ),
    .A2(_01849_),
    .B1(_01851_),
    .B2(\filters.cutoff_lut[9] ),
    .ZN(_01852_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09462_ (.I(_01827_),
    .Z(_01853_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09463_ (.A1(_00997_),
    .A2(_01784_),
    .ZN(_01854_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _09464_ (.A1(_01789_),
    .A2(_01853_),
    .A3(_01854_),
    .ZN(_01855_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09465_ (.A1(_00997_),
    .A2(net3),
    .ZN(_01856_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _09466_ (.A1(_01856_),
    .A2(_01789_),
    .A3(_01853_),
    .ZN(_01857_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09467_ (.A1(\channels.freq1[0] ),
    .A2(_01855_),
    .B1(_01857_),
    .B2(\channels.ctrl_reg1[0] ),
    .ZN(_01858_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09468_ (.A1(_01000_),
    .A2(_01789_),
    .ZN(_01859_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _09469_ (.A1(net2),
    .A2(_01787_),
    .A3(_01845_),
    .ZN(_01860_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09470_ (.A1(_01785_),
    .A2(_01860_),
    .ZN(_01861_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09471_ (.I(_01861_),
    .Z(_01862_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _09472_ (.A1(\channels.sus_rel3[0] ),
    .A2(_01859_),
    .B1(_01862_),
    .B2(\channels.pw2[8] ),
    .ZN(_01863_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _09473_ (.A1(_01852_),
    .A2(_01858_),
    .A3(_01863_),
    .ZN(_01864_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _09474_ (.A1(_01748_),
    .A2(_01844_),
    .B1(_01848_),
    .B2(\channels.pw2[0] ),
    .C(_01864_),
    .ZN(_01865_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09475_ (.A1(_01825_),
    .A2(_01840_),
    .ZN(_01866_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09476_ (.I(_01866_),
    .Z(_01867_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09477_ (.A1(_01832_),
    .A2(_01846_),
    .ZN(_01868_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09478_ (.I(_01868_),
    .Z(_01869_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09479_ (.A1(_01832_),
    .A2(_01860_),
    .ZN(_01870_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _09480_ (.I(_01870_),
    .Z(_01871_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_4 _09481_ (.A1(\channels.atk_dec3[0] ),
    .A2(_01867_),
    .B1(_01869_),
    .B2(\channels.sus_rel2[0] ),
    .C1(_01871_),
    .C2(\channels.freq3[0] ),
    .ZN(_01872_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _09482_ (.A1(_01835_),
    .A2(_01843_),
    .A3(_01865_),
    .A4(_01872_),
    .ZN(_01873_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09483_ (.I(net7),
    .Z(_01874_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09484_ (.I(_01874_),
    .Z(_01875_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _09485_ (.A1(_01783_),
    .A2(_01836_),
    .A3(_01831_),
    .ZN(_01876_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09486_ (.I(_01876_),
    .Z(_01877_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09487_ (.A1(\channels.ch3_env[0] ),
    .A2(_01877_),
    .ZN(_01878_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _09488_ (.A1(_01856_),
    .A2(_01824_),
    .A3(_01853_),
    .ZN(_01879_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09489_ (.I(_01879_),
    .Z(_01880_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09490_ (.A1(_01850_),
    .A2(_01840_),
    .ZN(_01881_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09491_ (.I(_01881_),
    .Z(_01882_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09492_ (.A1(\channels.freq2[0] ),
    .A2(_01880_),
    .B1(_01882_),
    .B2(\channels.ctrl_reg3[0] ),
    .ZN(_01883_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09493_ (.A1(_01854_),
    .A2(_01860_),
    .ZN(_01884_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09494_ (.I(_01884_),
    .Z(_01885_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09495_ (.A1(_01854_),
    .A2(_01846_),
    .ZN(_01886_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09496_ (.I(_01886_),
    .Z(_01887_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09497_ (.A1(\channels.pw1[0] ),
    .A2(_01885_),
    .B1(_01887_),
    .B2(\channels.freq1[8] ),
    .ZN(_01888_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _09498_ (.A1(_01875_),
    .A2(_01878_),
    .A3(_01883_),
    .A4(_01888_),
    .ZN(_01889_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _09499_ (.A1(_01825_),
    .A2(_01853_),
    .A3(_01854_),
    .ZN(_01890_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09500_ (.I(_01890_),
    .Z(_01891_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _09501_ (.A1(_01826_),
    .A2(_01836_),
    .A3(_01828_),
    .ZN(_01892_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09502_ (.I(_01892_),
    .Z(_01893_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09503_ (.A1(\channels.pw1[8] ),
    .A2(_01891_),
    .B1(_01893_),
    .B2(\channels.freq2[8] ),
    .ZN(_01894_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09504_ (.A1(_01836_),
    .A2(_01840_),
    .ZN(_01895_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09505_ (.I(_01895_),
    .Z(_01896_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09506_ (.A1(\filters.mode_vol[0] ),
    .A2(_01791_),
    .B1(_01896_),
    .B2(\channels.pw3[0] ),
    .ZN(_01897_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09507_ (.A1(_01856_),
    .A2(_01860_),
    .ZN(_01898_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09508_ (.I(_01898_),
    .Z(_01899_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09509_ (.A1(_01856_),
    .A2(_01846_),
    .ZN(_01900_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09510_ (.I(_01900_),
    .Z(_01901_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09511_ (.A1(\channels.sus_rel1[0] ),
    .A2(_01899_),
    .B1(_01901_),
    .B2(\channels.atk_dec1[0] ),
    .ZN(_01902_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _09512_ (.A1(_01783_),
    .A2(_01824_),
    .A3(_01785_),
    .ZN(_01903_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09513_ (.I(_01903_),
    .Z(_01904_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _09514_ (.A1(_01783_),
    .A2(_01826_),
    .A3(_01839_),
    .ZN(_01905_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09515_ (.A1(\channels.sample3[4] ),
    .A2(_01904_),
    .B1(_01905_),
    .B2(\clk_trg[0] ),
    .ZN(_01906_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _09516_ (.A1(_01894_),
    .A2(_01897_),
    .A3(_01902_),
    .A4(_01906_),
    .ZN(_01907_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09517_ (.I(_01874_),
    .Z(_01908_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09518_ (.I(_01908_),
    .Z(_01909_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _09519_ (.A1(_01873_),
    .A2(_01889_),
    .A3(_01907_),
    .B1(net22),
    .B2(_01909_),
    .ZN(_01910_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09520_ (.A1(_01823_),
    .A2(_01910_),
    .ZN(_00141_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _09521_ (.A1(\channels.ctrl_reg2[1] ),
    .A2(_01830_),
    .B1(_01834_),
    .B2(\channels.freq3[9] ),
    .ZN(_01911_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _09522_ (.A1(\channels.atk_dec2[1] ),
    .A2(_01838_),
    .B1(_01842_),
    .B2(\channels.pw3[9] ),
    .ZN(_01912_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _09523_ (.A1(\filters.cutoff_lut[7] ),
    .A2(_01849_),
    .B1(_01851_),
    .B2(\filters.cutoff_lut[10] ),
    .ZN(_01913_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09524_ (.A1(\channels.freq1[1] ),
    .A2(_01855_),
    .B1(_01857_),
    .B2(\channels.ctrl_reg1[1] ),
    .ZN(_01914_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _09525_ (.A1(\channels.sus_rel3[1] ),
    .A2(_01859_),
    .B1(_01861_),
    .B2(\channels.pw2[9] ),
    .ZN(_01915_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _09526_ (.A1(_01913_),
    .A2(_01914_),
    .A3(_01915_),
    .ZN(_01916_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _09527_ (.A1(_01762_),
    .A2(_01844_),
    .B1(_01848_),
    .B2(\channels.pw2[1] ),
    .C(_01916_),
    .ZN(_01917_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_4 _09528_ (.A1(\channels.atk_dec3[1] ),
    .A2(_01867_),
    .B1(_01869_),
    .B2(\channels.sus_rel2[1] ),
    .C1(_01871_),
    .C2(\channels.freq3[1] ),
    .ZN(_01918_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _09529_ (.A1(_01911_),
    .A2(_01912_),
    .A3(_01917_),
    .A4(_01918_),
    .ZN(_01919_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09530_ (.A1(\channels.ch3_env[1] ),
    .A2(_01877_),
    .ZN(_01920_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09531_ (.A1(\channels.freq2[1] ),
    .A2(_01880_),
    .B1(_01882_),
    .B2(\channels.ctrl_reg3[1] ),
    .ZN(_01921_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09532_ (.A1(\channels.pw1[1] ),
    .A2(_01885_),
    .B1(_01887_),
    .B2(\channels.freq1[9] ),
    .ZN(_01922_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _09533_ (.A1(_01875_),
    .A2(_01920_),
    .A3(_01921_),
    .A4(_01922_),
    .ZN(_01923_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09534_ (.A1(\channels.pw1[9] ),
    .A2(_01891_),
    .B1(_01893_),
    .B2(\channels.freq2[9] ),
    .ZN(_01924_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09535_ (.A1(\filters.mode_vol[1] ),
    .A2(_01791_),
    .B1(_01896_),
    .B2(\channels.pw3[1] ),
    .ZN(_01925_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09536_ (.A1(\channels.sus_rel1[1] ),
    .A2(_01899_),
    .B1(_01901_),
    .B2(\channels.atk_dec1[1] ),
    .ZN(_01926_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09537_ (.I(\channels.sample3[5] ),
    .Z(_01927_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09538_ (.A1(_01927_),
    .A2(_01904_),
    .B1(_01905_),
    .B2(\clk_trg[1] ),
    .ZN(_01928_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _09539_ (.A1(_01924_),
    .A2(_01925_),
    .A3(_01926_),
    .A4(_01928_),
    .ZN(_01929_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _09540_ (.A1(_01919_),
    .A2(_01923_),
    .A3(_01929_),
    .B1(net23),
    .B2(_01909_),
    .ZN(_01930_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09541_ (.A1(_01823_),
    .A2(_01930_),
    .ZN(_00142_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09542_ (.I(_01087_),
    .Z(_01931_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09543_ (.I(_01931_),
    .Z(_01932_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _09544_ (.I(_01932_),
    .Z(_01933_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09545_ (.I(_01874_),
    .Z(_01934_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09546_ (.A1(\channels.ctrl_reg3[2] ),
    .A2(_01882_),
    .B1(_01862_),
    .B2(\channels.pw2[10] ),
    .ZN(_01935_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09547_ (.I(_01868_),
    .Z(_01936_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09548_ (.I(_01870_),
    .Z(_01937_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09549_ (.A1(\channels.sus_rel2[2] ),
    .A2(_01936_),
    .B1(_01937_),
    .B2(\channels.freq3[2] ),
    .ZN(_01938_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09550_ (.I(_01904_),
    .Z(_01939_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09551_ (.A1(_01773_),
    .A2(_01002_),
    .B1(_01790_),
    .B2(\filters.mode_vol[2] ),
    .ZN(_01940_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09552_ (.I(_01857_),
    .Z(_01941_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09553_ (.A1(\channels.pw1[10] ),
    .A2(_01890_),
    .B1(_01941_),
    .B2(\channels.ctrl_reg1[2] ),
    .ZN(_01942_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09554_ (.I(_01859_),
    .Z(_01943_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09555_ (.A1(\filters.cutoff_lut[8] ),
    .A2(_01849_),
    .B1(_01943_),
    .B2(\channels.sus_rel3[2] ),
    .ZN(_01944_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09556_ (.A1(_01940_),
    .A2(_01942_),
    .A3(_01944_),
    .ZN(_01945_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _09557_ (.A1(\channels.sus_rel1[2] ),
    .A2(_01899_),
    .B1(_01939_),
    .B2(\channels.sample3[6] ),
    .C(_01945_),
    .ZN(_01946_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09558_ (.A1(_01935_),
    .A2(_01938_),
    .A3(_01946_),
    .ZN(_01947_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09559_ (.I(_01900_),
    .Z(_01948_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09560_ (.A1(\channels.atk_dec1[2] ),
    .A2(_01948_),
    .ZN(_01949_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09561_ (.A1(\channels.pw1[2] ),
    .A2(_01884_),
    .B1(_01892_),
    .B2(\channels.freq2[10] ),
    .ZN(_01950_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09562_ (.A1(\channels.ctrl_reg2[2] ),
    .A2(_01829_),
    .B1(_01879_),
    .B2(\channels.freq2[2] ),
    .ZN(_01951_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09563_ (.A1(_01950_),
    .A2(_01951_),
    .ZN(_01952_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _09564_ (.A1(\channels.pw3[10] ),
    .A2(_01842_),
    .B1(_01848_),
    .B2(\channels.pw2[2] ),
    .C(_01952_),
    .ZN(_01953_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09565_ (.I(_01855_),
    .Z(_01954_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09566_ (.A1(\channels.ch3_env[2] ),
    .A2(_01876_),
    .B1(_01886_),
    .B2(\channels.freq1[10] ),
    .ZN(_01955_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09567_ (.I(_01851_),
    .Z(_01956_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09568_ (.A1(\filters.cutoff_lut[11] ),
    .A2(_01956_),
    .B1(_01866_),
    .B2(\channels.atk_dec3[2] ),
    .ZN(_01957_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09569_ (.A1(\channels.atk_dec2[2] ),
    .A2(_01837_),
    .B1(_01895_),
    .B2(\channels.pw3[2] ),
    .ZN(_01958_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09570_ (.A1(_01955_),
    .A2(_01957_),
    .A3(_01958_),
    .ZN(_01959_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _09571_ (.A1(\channels.freq1[2] ),
    .A2(_01954_),
    .B1(_01834_),
    .B2(\channels.freq3[10] ),
    .C(_01959_),
    .ZN(_01960_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _09572_ (.A1(_01875_),
    .A2(_01949_),
    .A3(_01953_),
    .A4(_01960_),
    .ZN(_01961_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09573_ (.A1(_01934_),
    .A2(net24),
    .B1(_01947_),
    .B2(_01961_),
    .ZN(_01962_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09574_ (.A1(_01933_),
    .A2(_01962_),
    .ZN(_00143_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09575_ (.I(_01943_),
    .Z(_01963_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09576_ (.I(_01898_),
    .Z(_01964_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09577_ (.A1(\channels.sus_rel3[3] ),
    .A2(_01963_),
    .B1(_01964_),
    .B2(\channels.sus_rel1[3] ),
    .ZN(_01965_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09578_ (.I(_01837_),
    .Z(_01966_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09579_ (.A1(\filters.res_filt[3] ),
    .A2(_01844_),
    .B1(_01893_),
    .B2(\channels.freq2[11] ),
    .ZN(_01967_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09580_ (.A1(\filters.mode_vol[3] ),
    .A2(_01790_),
    .B1(_01868_),
    .B2(\channels.sus_rel2[3] ),
    .ZN(_01968_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09581_ (.A1(\channels.ch3_env[3] ),
    .A2(_01877_),
    .B1(_01885_),
    .B2(\channels.pw1[3] ),
    .ZN(_01969_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09582_ (.I(_01886_),
    .Z(_01970_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09583_ (.A1(\channels.pw3[11] ),
    .A2(_01841_),
    .B1(_01970_),
    .B2(\channels.freq1[11] ),
    .ZN(_01971_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _09584_ (.A1(_01967_),
    .A2(_01968_),
    .A3(_01969_),
    .A4(_01971_),
    .ZN(_01972_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09585_ (.A1(\channels.atk_dec2[3] ),
    .A2(_01966_),
    .B(_01972_),
    .ZN(_01973_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09586_ (.I(_01829_),
    .Z(_01974_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09587_ (.A1(\channels.pw1[11] ),
    .A2(_01891_),
    .ZN(_01975_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09588_ (.A1(\channels.freq3[3] ),
    .A2(_01870_),
    .B1(_01879_),
    .B2(\channels.freq2[3] ),
    .ZN(_01976_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09589_ (.I(\channels.sample3[7] ),
    .Z(_01977_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _09590_ (.A1(\channels.ctrl_reg1[3] ),
    .A2(_01941_),
    .B1(_01903_),
    .B2(_01977_),
    .ZN(_01978_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _09591_ (.A1(_01874_),
    .A2(_01975_),
    .A3(_01976_),
    .A4(_01978_),
    .ZN(_01979_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _09592_ (.A1(\channels.ctrl_reg2[3] ),
    .A2(_01974_),
    .B1(_01882_),
    .B2(\channels.ctrl_reg3[3] ),
    .C(_01979_),
    .ZN(_01980_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09593_ (.A1(\channels.pw2[3] ),
    .A2(_01847_),
    .B1(_01900_),
    .B2(\channels.atk_dec1[3] ),
    .ZN(_01981_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09594_ (.A1(\channels.atk_dec3[3] ),
    .A2(_01867_),
    .B1(_01895_),
    .B2(\channels.pw3[3] ),
    .ZN(_01982_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09595_ (.A1(\filters.cutoff_lut[12] ),
    .A2(_01956_),
    .B1(_01954_),
    .B2(\channels.freq1[3] ),
    .ZN(_01983_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09596_ (.A1(_01981_),
    .A2(_01982_),
    .A3(_01983_),
    .ZN(_01984_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _09597_ (.A1(\channels.freq3[11] ),
    .A2(_01834_),
    .B1(_01862_),
    .B2(\channels.pw2[11] ),
    .C(_01984_),
    .ZN(_01985_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _09598_ (.A1(_01965_),
    .A2(_01973_),
    .A3(_01980_),
    .A4(_01985_),
    .ZN(_01986_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09599_ (.A1(_01909_),
    .A2(net25),
    .B(_01986_),
    .ZN(_01987_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09600_ (.A1(_01933_),
    .A2(_01987_),
    .ZN(_00144_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09601_ (.I(_01956_),
    .Z(_01988_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09602_ (.A1(\filters.cutoff_lut[13] ),
    .A2(_01988_),
    .ZN(_01989_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09603_ (.A1(\channels.sus_rel3[4] ),
    .A2(_01963_),
    .B1(_01887_),
    .B2(\channels.freq1[12] ),
    .ZN(_01990_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09604_ (.I(_01866_),
    .Z(_01991_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09605_ (.I(_01833_),
    .Z(_01992_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _09606_ (.A1(\channels.atk_dec3[4] ),
    .A2(_01991_),
    .B1(_01992_),
    .B2(\channels.freq3[12] ),
    .ZN(_01993_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _09607_ (.A1(_01875_),
    .A2(_01989_),
    .A3(_01990_),
    .A4(_01993_),
    .ZN(_01994_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _09608_ (.A1(\channels.ctrl_reg2[4] ),
    .A2(_01974_),
    .B1(_01966_),
    .B2(\channels.atk_dec2[4] ),
    .C(_01994_),
    .ZN(_01995_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09609_ (.I(_01847_),
    .Z(_01996_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09610_ (.I(_01892_),
    .Z(_01997_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09611_ (.A1(\channels.pw2[4] ),
    .A2(_01996_),
    .B1(_01997_),
    .B2(\channels.freq2[12] ),
    .ZN(_01998_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09612_ (.I(_01881_),
    .Z(_01999_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09613_ (.A1(\channels.freq3[4] ),
    .A2(_01937_),
    .B1(_01999_),
    .B2(\channels.ctrl_reg3[4] ),
    .ZN(_02000_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09614_ (.I(_01880_),
    .Z(_02001_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09615_ (.A1(\channels.sus_rel2[4] ),
    .A2(_01936_),
    .B1(_02001_),
    .B2(\channels.freq2[4] ),
    .ZN(_02002_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09616_ (.I(_01884_),
    .Z(_02003_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09617_ (.I(_01941_),
    .Z(_02004_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09618_ (.A1(\channels.pw1[4] ),
    .A2(_02003_),
    .B1(_02004_),
    .B2(\channels.ctrl_reg1[4] ),
    .ZN(_02005_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _09619_ (.A1(_01998_),
    .A2(_02000_),
    .A3(_02002_),
    .A4(_02005_),
    .ZN(_02006_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09620_ (.I(_01844_),
    .Z(_02007_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _09621_ (.A1(\filters.res_filt[4] ),
    .A2(_02007_),
    .B1(_01939_),
    .B2(\channels.sample3[8] ),
    .ZN(_02008_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09622_ (.I(_01877_),
    .Z(_02009_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09623_ (.A1(\channels.ch3_env[4] ),
    .A2(_02009_),
    .B1(_01948_),
    .B2(\channels.atk_dec1[4] ),
    .ZN(_02010_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09624_ (.I(_01954_),
    .Z(_02011_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09625_ (.I(_01896_),
    .Z(_02012_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09626_ (.A1(\channels.freq1[4] ),
    .A2(_02011_),
    .B1(_02012_),
    .B2(\channels.pw3[4] ),
    .ZN(_02013_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09627_ (.I(_01791_),
    .Z(_02014_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09628_ (.A1(\filters.lp ),
    .A2(_02014_),
    .B1(_01964_),
    .B2(\channels.sus_rel1[4] ),
    .ZN(_02015_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _09629_ (.A1(_02008_),
    .A2(_02010_),
    .A3(_02013_),
    .A4(_02015_),
    .ZN(_02016_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09630_ (.A1(_02006_),
    .A2(_02016_),
    .ZN(_02017_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09631_ (.A1(_01934_),
    .A2(net26),
    .B(_01809_),
    .ZN(_02018_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09632_ (.A1(_01995_),
    .A2(_02017_),
    .B(_02018_),
    .ZN(_00145_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09633_ (.A1(\filters.cutoff_lut[14] ),
    .A2(_01988_),
    .ZN(_02019_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09634_ (.A1(\channels.sus_rel3[5] ),
    .A2(_01963_),
    .B1(_01970_),
    .B2(\channels.freq1[13] ),
    .ZN(_02020_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _09635_ (.A1(\channels.atk_dec3[5] ),
    .A2(_01991_),
    .B1(_01992_),
    .B2(\channels.freq3[13] ),
    .ZN(_02021_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _09636_ (.A1(_01908_),
    .A2(_02019_),
    .A3(_02020_),
    .A4(_02021_),
    .ZN(_02022_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _09637_ (.A1(\channels.ctrl_reg2[5] ),
    .A2(_01974_),
    .B1(_01966_),
    .B2(\channels.atk_dec2[5] ),
    .C(_02022_),
    .ZN(_02023_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09638_ (.A1(\channels.pw2[5] ),
    .A2(_01996_),
    .B1(_01997_),
    .B2(\channels.freq2[13] ),
    .ZN(_02024_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09639_ (.A1(\channels.freq3[5] ),
    .A2(_01937_),
    .B1(_01999_),
    .B2(\channels.ctrl_reg3[5] ),
    .ZN(_02025_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09640_ (.A1(\channels.sus_rel2[5] ),
    .A2(_01936_),
    .B1(_02001_),
    .B2(\channels.freq2[5] ),
    .ZN(_02026_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09641_ (.A1(\channels.pw1[5] ),
    .A2(_02003_),
    .B1(_02004_),
    .B2(\channels.ctrl_reg1[5] ),
    .ZN(_02027_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _09642_ (.A1(_02024_),
    .A2(_02025_),
    .A3(_02026_),
    .A4(_02027_),
    .ZN(_02028_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09643_ (.I(\channels.sample3[9] ),
    .Z(_02029_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _09644_ (.A1(\filters.res_filt[5] ),
    .A2(_02007_),
    .B1(_01939_),
    .B2(_02029_),
    .ZN(_02030_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09645_ (.A1(\channels.ch3_env[5] ),
    .A2(_02009_),
    .B1(_01948_),
    .B2(\channels.atk_dec1[5] ),
    .ZN(_02031_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09646_ (.A1(\channels.freq1[5] ),
    .A2(_02011_),
    .B1(_02012_),
    .B2(\channels.pw3[5] ),
    .ZN(_02032_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _09647_ (.A1(\filters.bp ),
    .A2(_02014_),
    .B1(_01964_),
    .B2(\channels.sus_rel1[5] ),
    .ZN(_02033_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _09648_ (.A1(_02030_),
    .A2(_02031_),
    .A3(_02032_),
    .A4(_02033_),
    .ZN(_02034_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09649_ (.A1(_02028_),
    .A2(_02034_),
    .ZN(_02035_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09650_ (.I(_01808_),
    .Z(_02036_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09651_ (.A1(_01934_),
    .A2(net27),
    .B(_02036_),
    .ZN(_02037_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09652_ (.A1(_02023_),
    .A2(_02035_),
    .B(_02037_),
    .ZN(_00146_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09653_ (.A1(\filters.cutoff_lut[15] ),
    .A2(_01988_),
    .ZN(_02038_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09654_ (.A1(\channels.sus_rel3[6] ),
    .A2(_01943_),
    .B1(_01970_),
    .B2(\channels.freq1[14] ),
    .ZN(_02039_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09655_ (.A1(\channels.atk_dec3[6] ),
    .A2(_01991_),
    .B1(_01992_),
    .B2(\channels.freq3[14] ),
    .ZN(_02040_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _09656_ (.A1(_01908_),
    .A2(_02038_),
    .A3(_02039_),
    .A4(_02040_),
    .ZN(_02041_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _09657_ (.A1(\channels.ctrl_reg2[6] ),
    .A2(_01974_),
    .B1(_01966_),
    .B2(\channels.atk_dec2[6] ),
    .C(_02041_),
    .ZN(_02042_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09658_ (.A1(\channels.pw2[6] ),
    .A2(_01996_),
    .B1(_01997_),
    .B2(\channels.freq2[14] ),
    .ZN(_02043_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09659_ (.A1(\channels.freq3[6] ),
    .A2(_01871_),
    .B1(_01999_),
    .B2(\channels.ctrl_reg3[6] ),
    .ZN(_02044_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09660_ (.A1(\channels.sus_rel2[6] ),
    .A2(_01869_),
    .B1(_02001_),
    .B2(\channels.freq2[6] ),
    .ZN(_02045_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09661_ (.A1(\channels.pw1[6] ),
    .A2(_02003_),
    .B1(_02004_),
    .B2(\channels.ctrl_reg1[6] ),
    .ZN(_02046_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _09662_ (.A1(_02043_),
    .A2(_02044_),
    .A3(_02045_),
    .A4(_02046_),
    .ZN(_02047_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _09663_ (.A1(\filters.res_filt[6] ),
    .A2(_02007_),
    .B1(_01939_),
    .B2(\channels.sample3[10] ),
    .ZN(_02048_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09664_ (.A1(\channels.ch3_env[6] ),
    .A2(_02009_),
    .B1(_01948_),
    .B2(\channels.atk_dec1[6] ),
    .ZN(_02049_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09665_ (.A1(\channels.freq1[6] ),
    .A2(_02011_),
    .B1(_02012_),
    .B2(\channels.pw3[6] ),
    .ZN(_02050_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09666_ (.A1(\filters.hp ),
    .A2(_02014_),
    .B1(_01899_),
    .B2(\channels.sus_rel1[6] ),
    .ZN(_02051_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _09667_ (.A1(_02048_),
    .A2(_02049_),
    .A3(_02050_),
    .A4(_02051_),
    .ZN(_02052_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09668_ (.A1(_02047_),
    .A2(_02052_),
    .ZN(_02053_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09669_ (.A1(_01934_),
    .A2(net28),
    .B(_02036_),
    .ZN(_02054_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09670_ (.A1(_02042_),
    .A2(_02053_),
    .B(_02054_),
    .ZN(_00147_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _09671_ (.A1(\channels.atk_dec3[7] ),
    .A2(_01991_),
    .B1(_01992_),
    .B2(\channels.freq3[15] ),
    .ZN(_02055_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09672_ (.I(\channels.sample3[11] ),
    .Z(_02056_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09673_ (.A1(\channels.ctrl_reg2[7] ),
    .A2(_01830_),
    .B1(_01904_),
    .B2(_02056_),
    .ZN(_02057_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09674_ (.A1(\channels.atk_dec1[7] ),
    .A2(_01901_),
    .B(_01905_),
    .ZN(_02058_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _09675_ (.A1(_01908_),
    .A2(_02055_),
    .A3(_02057_),
    .A4(_02058_),
    .ZN(_02059_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _09676_ (.A1(\channels.sus_rel3[7] ),
    .A2(_01963_),
    .B1(_01964_),
    .B2(\channels.sus_rel1[7] ),
    .C(_02059_),
    .ZN(_02060_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09677_ (.A1(\channels.freq1[7] ),
    .A2(_02011_),
    .B1(_01936_),
    .B2(\channels.sus_rel2[7] ),
    .ZN(_02061_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09678_ (.A1(\filters.mode_vol[7] ),
    .A2(_02014_),
    .B1(_02001_),
    .B2(\channels.freq2[7] ),
    .ZN(_02062_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09679_ (.A1(\channels.freq2[15] ),
    .A2(_01997_),
    .B1(_01887_),
    .B2(\channels.freq1[15] ),
    .ZN(_02063_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09680_ (.A1(\channels.atk_dec2[7] ),
    .A2(_01838_),
    .B1(_01937_),
    .B2(\channels.freq3[7] ),
    .ZN(_02064_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _09681_ (.A1(_02061_),
    .A2(_02062_),
    .A3(_02063_),
    .A4(_02064_),
    .ZN(_02065_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09682_ (.A1(\channels.ctrl_reg3[7] ),
    .A2(_01999_),
    .B1(_02004_),
    .B2(\channels.ctrl_reg1[7] ),
    .ZN(_02066_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09683_ (.A1(\filters.cutoff_lut[16] ),
    .A2(_01988_),
    .B1(_02009_),
    .B2(\channels.ch3_env[7] ),
    .ZN(_02067_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09684_ (.A1(\filters.res_filt[7] ),
    .A2(_02007_),
    .B1(_02012_),
    .B2(\channels.pw3[7] ),
    .ZN(_02068_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09685_ (.A1(\channels.pw1[7] ),
    .A2(_02003_),
    .B1(_01996_),
    .B2(\channels.pw2[7] ),
    .ZN(_02069_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _09686_ (.A1(_02066_),
    .A2(_02067_),
    .A3(_02068_),
    .A4(_02069_),
    .ZN(_02070_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09687_ (.A1(_02065_),
    .A2(_02070_),
    .ZN(_02071_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09688_ (.A1(net29),
    .A2(_01909_),
    .B(_02036_),
    .ZN(_02072_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09689_ (.A1(_02060_),
    .A2(_02071_),
    .B(_02072_),
    .ZN(_00148_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09690_ (.A1(_01781_),
    .A2(_01970_),
    .Z(_02073_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09691_ (.I(_02073_),
    .Z(_02074_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09692_ (.I(_02073_),
    .Z(_02075_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09693_ (.A1(\channels.freq1[8] ),
    .A2(_02075_),
    .B(_02036_),
    .ZN(_02076_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09694_ (.A1(_01742_),
    .A2(_02074_),
    .B(_02076_),
    .ZN(_00149_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09695_ (.I(_01808_),
    .Z(_02077_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09696_ (.A1(\channels.freq1[9] ),
    .A2(_02075_),
    .B(_02077_),
    .ZN(_02078_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09697_ (.A1(_01757_),
    .A2(_02074_),
    .B(_02078_),
    .ZN(_00150_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09698_ (.A1(\channels.freq1[10] ),
    .A2(_02075_),
    .B(_02077_),
    .ZN(_02079_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09699_ (.A1(_01767_),
    .A2(_02074_),
    .B(_02079_),
    .ZN(_00151_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09700_ (.A1(\channels.freq1[11] ),
    .A2(_02075_),
    .B(_02077_),
    .ZN(_02080_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09701_ (.A1(_01777_),
    .A2(_02074_),
    .B(_02080_),
    .ZN(_00152_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09702_ (.I(_02073_),
    .Z(_02081_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09703_ (.I(_02073_),
    .Z(_02082_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09704_ (.A1(\channels.freq1[12] ),
    .A2(_02082_),
    .B(_02077_),
    .ZN(_02083_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09705_ (.A1(_01801_),
    .A2(_02081_),
    .B(_02083_),
    .ZN(_00153_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09706_ (.I(_01808_),
    .Z(_02084_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09707_ (.A1(\channels.freq1[13] ),
    .A2(_02082_),
    .B(_02084_),
    .ZN(_02085_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09708_ (.A1(_01807_),
    .A2(_02081_),
    .B(_02085_),
    .ZN(_00154_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09709_ (.A1(\channels.freq1[14] ),
    .A2(_02082_),
    .B(_02084_),
    .ZN(_02086_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09710_ (.A1(_01814_),
    .A2(_02081_),
    .B(_02086_),
    .ZN(_00155_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09711_ (.A1(\channels.freq1[15] ),
    .A2(_02082_),
    .B(_02084_),
    .ZN(_02087_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09712_ (.A1(_01819_),
    .A2(_02081_),
    .B(_02087_),
    .ZN(_00156_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09713_ (.I(_01780_),
    .Z(_02088_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09714_ (.A1(_02088_),
    .A2(_01891_),
    .Z(_02089_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09715_ (.I(_02089_),
    .Z(_02090_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09716_ (.I(_02089_),
    .Z(_02091_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09717_ (.A1(\channels.pw1[8] ),
    .A2(_02091_),
    .B(_02084_),
    .ZN(_02092_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09718_ (.A1(_01742_),
    .A2(_02090_),
    .B(_02092_),
    .ZN(_00157_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09719_ (.I(_01751_),
    .Z(_02093_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09720_ (.I(_02093_),
    .Z(_02094_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09721_ (.A1(\channels.pw1[9] ),
    .A2(_02091_),
    .B(_02094_),
    .ZN(_02095_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09722_ (.A1(_01757_),
    .A2(_02090_),
    .B(_02095_),
    .ZN(_00158_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09723_ (.A1(\channels.pw1[10] ),
    .A2(_02091_),
    .B(_02094_),
    .ZN(_02096_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09724_ (.A1(_01767_),
    .A2(_02090_),
    .B(_02096_),
    .ZN(_00159_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09725_ (.I(\channels.pw1[11] ),
    .ZN(_02097_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09726_ (.I(net11),
    .Z(_02098_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09727_ (.A1(_02098_),
    .A2(_02091_),
    .ZN(_02099_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09728_ (.I(_01062_),
    .Z(_02100_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09729_ (.I(_02100_),
    .Z(_02101_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09730_ (.I(_02101_),
    .Z(_02102_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09731_ (.I(_02102_),
    .Z(_02103_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09732_ (.A1(_02097_),
    .A2(_02090_),
    .B(_02099_),
    .C(_02103_),
    .ZN(_00160_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09733_ (.I(_01739_),
    .Z(_02104_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09734_ (.I(_02104_),
    .Z(_02105_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09735_ (.A1(_01781_),
    .A2(_01941_),
    .Z(_02106_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09736_ (.I(_02106_),
    .Z(_02107_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09737_ (.I(_02106_),
    .Z(_02108_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09738_ (.A1(\channels.ctrl_reg1[0] ),
    .A2(_02108_),
    .B(_02094_),
    .ZN(_02109_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09739_ (.A1(_02105_),
    .A2(_02107_),
    .B(_02109_),
    .ZN(_00161_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09740_ (.I(_01756_),
    .Z(_02110_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09741_ (.A1(\channels.ctrl_reg1[1] ),
    .A2(_02108_),
    .B(_02094_),
    .ZN(_02111_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09742_ (.A1(_02110_),
    .A2(_02107_),
    .B(_02111_),
    .ZN(_00162_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09743_ (.I(_01766_),
    .Z(_02112_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09744_ (.I(_02093_),
    .Z(_02113_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09745_ (.A1(\channels.ctrl_reg1[2] ),
    .A2(_02108_),
    .B(_02113_),
    .ZN(_02114_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09746_ (.A1(_02112_),
    .A2(_02107_),
    .B(_02114_),
    .ZN(_00163_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09747_ (.A1(\channels.ctrl_reg1[3] ),
    .A2(_02108_),
    .B(_02113_),
    .ZN(_02115_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09748_ (.A1(_01777_),
    .A2(_02107_),
    .B(_02115_),
    .ZN(_00164_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09749_ (.I(_02106_),
    .Z(_02116_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09750_ (.I(_02106_),
    .Z(_02117_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09751_ (.A1(\channels.ctrl_reg1[4] ),
    .A2(_02117_),
    .B(_02113_),
    .ZN(_02118_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09752_ (.A1(_01801_),
    .A2(_02116_),
    .B(_02118_),
    .ZN(_00165_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09753_ (.A1(\channels.ctrl_reg1[5] ),
    .A2(_02117_),
    .B(_02113_),
    .ZN(_02119_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09754_ (.A1(_01807_),
    .A2(_02116_),
    .B(_02119_),
    .ZN(_00166_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09755_ (.I(_02093_),
    .Z(_02120_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09756_ (.A1(\channels.ctrl_reg1[6] ),
    .A2(_02117_),
    .B(_02120_),
    .ZN(_02121_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09757_ (.A1(_01814_),
    .A2(_02116_),
    .B(_02121_),
    .ZN(_00167_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09758_ (.A1(\channels.ctrl_reg1[7] ),
    .A2(_02117_),
    .B(_02120_),
    .ZN(_02122_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09759_ (.A1(_01819_),
    .A2(_02116_),
    .B(_02122_),
    .ZN(_00168_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09760_ (.I(_01780_),
    .Z(_02123_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09761_ (.A1(_02123_),
    .A2(_01901_),
    .Z(_02124_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09762_ (.I(_02124_),
    .Z(_02125_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09763_ (.I(_02124_),
    .Z(_02126_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09764_ (.A1(\channels.atk_dec1[0] ),
    .A2(_02126_),
    .B(_02120_),
    .ZN(_02127_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09765_ (.A1(_02105_),
    .A2(_02125_),
    .B(_02127_),
    .ZN(_00169_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09766_ (.A1(\channels.atk_dec1[1] ),
    .A2(_02126_),
    .B(_02120_),
    .ZN(_02128_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09767_ (.A1(_02110_),
    .A2(_02125_),
    .B(_02128_),
    .ZN(_00170_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09768_ (.I(_02093_),
    .Z(_02129_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09769_ (.A1(\channels.atk_dec1[2] ),
    .A2(_02126_),
    .B(_02129_),
    .ZN(_02130_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09770_ (.A1(_02112_),
    .A2(_02125_),
    .B(_02130_),
    .ZN(_00171_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09771_ (.I(_01776_),
    .Z(_02131_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09772_ (.A1(\channels.atk_dec1[3] ),
    .A2(_02126_),
    .B(_02129_),
    .ZN(_02132_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09773_ (.A1(_02131_),
    .A2(_02125_),
    .B(_02132_),
    .ZN(_00172_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09774_ (.I(_02124_),
    .Z(_02133_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09775_ (.I(_02124_),
    .Z(_02134_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09776_ (.A1(\channels.atk_dec1[4] ),
    .A2(_02134_),
    .B(_02129_),
    .ZN(_02135_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09777_ (.A1(_01801_),
    .A2(_02133_),
    .B(_02135_),
    .ZN(_00173_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09778_ (.A1(\channels.atk_dec1[5] ),
    .A2(_02134_),
    .B(_02129_),
    .ZN(_02136_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09779_ (.A1(_01807_),
    .A2(_02133_),
    .B(_02136_),
    .ZN(_00174_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09780_ (.I(_01751_),
    .Z(_02137_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09781_ (.I(_02137_),
    .Z(_02138_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09782_ (.A1(\channels.atk_dec1[6] ),
    .A2(_02134_),
    .B(_02138_),
    .ZN(_02139_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09783_ (.A1(_01814_),
    .A2(_02133_),
    .B(_02139_),
    .ZN(_00175_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09784_ (.A1(\channels.atk_dec1[7] ),
    .A2(_02134_),
    .B(_02138_),
    .ZN(_02140_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09785_ (.A1(_01819_),
    .A2(_02133_),
    .B(_02140_),
    .ZN(_00176_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09786_ (.A1(_02123_),
    .A2(_01898_),
    .Z(_02141_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09787_ (.I(_02141_),
    .Z(_02142_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09788_ (.I(_02141_),
    .Z(_02143_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09789_ (.A1(\channels.sus_rel1[0] ),
    .A2(_02143_),
    .B(_02138_),
    .ZN(_02144_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09790_ (.A1(_02105_),
    .A2(_02142_),
    .B(_02144_),
    .ZN(_00177_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09791_ (.A1(\channels.sus_rel1[1] ),
    .A2(_02143_),
    .B(_02138_),
    .ZN(_02145_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09792_ (.A1(_02110_),
    .A2(_02142_),
    .B(_02145_),
    .ZN(_00178_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09793_ (.I(_02137_),
    .Z(_02146_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09794_ (.A1(\channels.sus_rel1[2] ),
    .A2(_02143_),
    .B(_02146_),
    .ZN(_02147_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09795_ (.A1(_02112_),
    .A2(_02142_),
    .B(_02147_),
    .ZN(_00179_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09796_ (.A1(\channels.sus_rel1[3] ),
    .A2(_02143_),
    .B(_02146_),
    .ZN(_02148_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09797_ (.A1(_02131_),
    .A2(_02142_),
    .B(_02148_),
    .ZN(_00180_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09798_ (.I(_01017_),
    .Z(_02149_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09799_ (.I(_02149_),
    .Z(_02150_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09800_ (.I(_02141_),
    .Z(_02151_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09801_ (.I(_02141_),
    .Z(_02152_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09802_ (.A1(\channels.sus_rel1[4] ),
    .A2(_02152_),
    .B(_02146_),
    .ZN(_02153_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09803_ (.A1(_02150_),
    .A2(_02151_),
    .B(_02153_),
    .ZN(_00181_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09804_ (.I(_01805_),
    .Z(_02154_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09805_ (.I(_02154_),
    .Z(_02155_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09806_ (.A1(\channels.sus_rel1[5] ),
    .A2(_02152_),
    .B(_02146_),
    .ZN(_02156_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09807_ (.A1(_02155_),
    .A2(_02151_),
    .B(_02156_),
    .ZN(_00182_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09808_ (.I(_01813_),
    .Z(_02157_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09809_ (.I(_02137_),
    .Z(_02158_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09810_ (.A1(\channels.sus_rel1[6] ),
    .A2(_02152_),
    .B(_02158_),
    .ZN(_02159_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09811_ (.A1(_02157_),
    .A2(_02151_),
    .B(_02159_),
    .ZN(_00183_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09812_ (.I(_01818_),
    .Z(_02160_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09813_ (.A1(\channels.sus_rel1[7] ),
    .A2(_02152_),
    .B(_02158_),
    .ZN(_02161_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09814_ (.A1(_02160_),
    .A2(_02151_),
    .B(_02161_),
    .ZN(_00184_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09815_ (.A1(_02123_),
    .A2(_01893_),
    .Z(_02162_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09816_ (.I(_02162_),
    .Z(_02163_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09817_ (.I(_02162_),
    .Z(_02164_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09818_ (.A1(\channels.freq2[8] ),
    .A2(_02164_),
    .B(_02158_),
    .ZN(_02165_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09819_ (.A1(_02105_),
    .A2(_02163_),
    .B(_02165_),
    .ZN(_00185_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09820_ (.A1(\channels.freq2[9] ),
    .A2(_02164_),
    .B(_02158_),
    .ZN(_02166_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09821_ (.A1(_02110_),
    .A2(_02163_),
    .B(_02166_),
    .ZN(_00186_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09822_ (.I(_02137_),
    .Z(_02167_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09823_ (.A1(\channels.freq2[10] ),
    .A2(_02164_),
    .B(_02167_),
    .ZN(_02168_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09824_ (.A1(_02112_),
    .A2(_02163_),
    .B(_02168_),
    .ZN(_00187_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09825_ (.A1(\channels.freq2[11] ),
    .A2(_02164_),
    .B(_02167_),
    .ZN(_02169_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09826_ (.A1(_02131_),
    .A2(_02163_),
    .B(_02169_),
    .ZN(_00188_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09827_ (.I(_02162_),
    .Z(_02170_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09828_ (.I(_02162_),
    .Z(_02171_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09829_ (.A1(\channels.freq2[12] ),
    .A2(_02171_),
    .B(_02167_),
    .ZN(_02172_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09830_ (.A1(_02150_),
    .A2(_02170_),
    .B(_02172_),
    .ZN(_00189_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09831_ (.A1(\channels.freq2[13] ),
    .A2(_02171_),
    .B(_02167_),
    .ZN(_02173_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09832_ (.A1(_02155_),
    .A2(_02170_),
    .B(_02173_),
    .ZN(_00190_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09833_ (.I(_01750_),
    .Z(_02174_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09834_ (.I(_02174_),
    .Z(_02175_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09835_ (.I(_02175_),
    .Z(_02176_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09836_ (.A1(\channels.freq2[14] ),
    .A2(_02171_),
    .B(_02176_),
    .ZN(_02177_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09837_ (.A1(_02157_),
    .A2(_02170_),
    .B(_02177_),
    .ZN(_00191_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09838_ (.A1(\channels.freq2[15] ),
    .A2(_02171_),
    .B(_02176_),
    .ZN(_02178_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09839_ (.A1(_02160_),
    .A2(_02170_),
    .B(_02178_),
    .ZN(_00192_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09840_ (.I(_02104_),
    .Z(_02179_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09841_ (.A1(_02088_),
    .A2(_01862_),
    .Z(_02180_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09842_ (.I(_02180_),
    .Z(_02181_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09843_ (.I(_02180_),
    .Z(_02182_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09844_ (.A1(\channels.pw2[8] ),
    .A2(_02182_),
    .B(_02176_),
    .ZN(_02183_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09845_ (.A1(_02179_),
    .A2(_02181_),
    .B(_02183_),
    .ZN(_00193_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09846_ (.I(_01755_),
    .Z(_02184_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09847_ (.I(_02184_),
    .Z(_02185_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09848_ (.A1(\channels.pw2[9] ),
    .A2(_02182_),
    .B(_02176_),
    .ZN(_02186_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09849_ (.A1(_02185_),
    .A2(_02181_),
    .B(_02186_),
    .ZN(_00194_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09850_ (.I(_01765_),
    .Z(_02187_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09851_ (.I(_02187_),
    .Z(_02188_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09852_ (.I(_02175_),
    .Z(_02189_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09853_ (.A1(\channels.pw2[10] ),
    .A2(_02182_),
    .B(_02189_),
    .ZN(_02190_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09854_ (.A1(_02188_),
    .A2(_02181_),
    .B(_02190_),
    .ZN(_00195_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09855_ (.I(\channels.pw2[11] ),
    .ZN(_02191_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09856_ (.A1(_02098_),
    .A2(_02182_),
    .ZN(_02192_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09857_ (.A1(_02191_),
    .A2(_02181_),
    .B(_02192_),
    .C(_02103_),
    .ZN(_00196_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09858_ (.A1(_02123_),
    .A2(_01830_),
    .Z(_02193_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09859_ (.I(_02193_),
    .Z(_02194_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09860_ (.I(_02193_),
    .Z(_02195_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09861_ (.A1(\channels.ctrl_reg2[0] ),
    .A2(_02195_),
    .B(_02189_),
    .ZN(_02196_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09862_ (.A1(_02179_),
    .A2(_02194_),
    .B(_02196_),
    .ZN(_00197_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09863_ (.A1(\channels.ctrl_reg2[1] ),
    .A2(_02195_),
    .B(_02189_),
    .ZN(_02197_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09864_ (.A1(_02185_),
    .A2(_02194_),
    .B(_02197_),
    .ZN(_00198_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09865_ (.A1(\channels.ctrl_reg2[2] ),
    .A2(_02195_),
    .B(_02189_),
    .ZN(_02198_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09866_ (.A1(_02188_),
    .A2(_02194_),
    .B(_02198_),
    .ZN(_00199_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09867_ (.I(_02175_),
    .Z(_02199_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09868_ (.A1(\channels.ctrl_reg2[3] ),
    .A2(_02195_),
    .B(_02199_),
    .ZN(_02200_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09869_ (.A1(_02131_),
    .A2(_02194_),
    .B(_02200_),
    .ZN(_00200_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09870_ (.I(_02193_),
    .Z(_02201_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09871_ (.I(_02193_),
    .Z(_02202_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09872_ (.A1(\channels.ctrl_reg2[4] ),
    .A2(_02202_),
    .B(_02199_),
    .ZN(_02203_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09873_ (.A1(_02150_),
    .A2(_02201_),
    .B(_02203_),
    .ZN(_00201_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09874_ (.A1(\channels.ctrl_reg2[5] ),
    .A2(_02202_),
    .B(_02199_),
    .ZN(_02204_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09875_ (.A1(_02155_),
    .A2(_02201_),
    .B(_02204_),
    .ZN(_00202_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09876_ (.A1(\channels.ctrl_reg2[6] ),
    .A2(_02202_),
    .B(_02199_),
    .ZN(_02205_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09877_ (.A1(_02157_),
    .A2(_02201_),
    .B(_02205_),
    .ZN(_00203_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09878_ (.I(_02175_),
    .Z(_02206_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09879_ (.A1(\channels.ctrl_reg2[7] ),
    .A2(_02202_),
    .B(_02206_),
    .ZN(_02207_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09880_ (.A1(_02160_),
    .A2(_02201_),
    .B(_02207_),
    .ZN(_00204_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09881_ (.I(_01779_),
    .Z(_02208_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09882_ (.A1(_02208_),
    .A2(_01838_),
    .Z(_02209_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09883_ (.I(_02209_),
    .Z(_02210_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09884_ (.I(_02209_),
    .Z(_02211_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09885_ (.A1(\channels.atk_dec2[0] ),
    .A2(_02211_),
    .B(_02206_),
    .ZN(_02212_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09886_ (.A1(_02179_),
    .A2(_02210_),
    .B(_02212_),
    .ZN(_00205_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09887_ (.A1(\channels.atk_dec2[1] ),
    .A2(_02211_),
    .B(_02206_),
    .ZN(_02213_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09888_ (.A1(_02185_),
    .A2(_02210_),
    .B(_02213_),
    .ZN(_00206_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09889_ (.A1(\channels.atk_dec2[2] ),
    .A2(_02211_),
    .B(_02206_),
    .ZN(_02214_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09890_ (.A1(_02188_),
    .A2(_02210_),
    .B(_02214_),
    .ZN(_00207_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09891_ (.I(_01776_),
    .Z(_02215_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09892_ (.I(_02174_),
    .Z(_02216_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09893_ (.I(_02216_),
    .Z(_02217_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09894_ (.A1(\channels.atk_dec2[3] ),
    .A2(_02211_),
    .B(_02217_),
    .ZN(_02218_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09895_ (.A1(_02215_),
    .A2(_02210_),
    .B(_02218_),
    .ZN(_00208_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09896_ (.I(_02209_),
    .Z(_02219_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09897_ (.I(_02209_),
    .Z(_02220_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09898_ (.A1(\channels.atk_dec2[4] ),
    .A2(_02220_),
    .B(_02217_),
    .ZN(_02221_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09899_ (.A1(_02150_),
    .A2(_02219_),
    .B(_02221_),
    .ZN(_00209_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09900_ (.A1(\channels.atk_dec2[5] ),
    .A2(_02220_),
    .B(_02217_),
    .ZN(_02222_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09901_ (.A1(_02155_),
    .A2(_02219_),
    .B(_02222_),
    .ZN(_00210_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09902_ (.A1(\channels.atk_dec2[6] ),
    .A2(_02220_),
    .B(_02217_),
    .ZN(_02223_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09903_ (.A1(_02157_),
    .A2(_02219_),
    .B(_02223_),
    .ZN(_00211_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09904_ (.I(_02216_),
    .Z(_02224_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09905_ (.A1(\channels.atk_dec2[7] ),
    .A2(_02220_),
    .B(_02224_),
    .ZN(_02225_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09906_ (.A1(_02160_),
    .A2(_02219_),
    .B(_02225_),
    .ZN(_00212_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09907_ (.A1(_02208_),
    .A2(_01869_),
    .Z(_02226_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09908_ (.I(_02226_),
    .Z(_02227_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09909_ (.I(_02226_),
    .Z(_02228_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09910_ (.A1(\channels.sus_rel2[0] ),
    .A2(_02228_),
    .B(_02224_),
    .ZN(_02229_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09911_ (.A1(_02179_),
    .A2(_02227_),
    .B(_02229_),
    .ZN(_00213_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09912_ (.A1(\channels.sus_rel2[1] ),
    .A2(_02228_),
    .B(_02224_),
    .ZN(_02230_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09913_ (.A1(_02185_),
    .A2(_02227_),
    .B(_02230_),
    .ZN(_00214_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09914_ (.A1(\channels.sus_rel2[2] ),
    .A2(_02228_),
    .B(_02224_),
    .ZN(_02231_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09915_ (.A1(_02188_),
    .A2(_02227_),
    .B(_02231_),
    .ZN(_00215_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09916_ (.I(_02216_),
    .Z(_02232_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09917_ (.A1(\channels.sus_rel2[3] ),
    .A2(_02228_),
    .B(_02232_),
    .ZN(_02233_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09918_ (.A1(_02215_),
    .A2(_02227_),
    .B(_02233_),
    .ZN(_00216_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09919_ (.I(_02149_),
    .Z(_02234_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09920_ (.I(_02226_),
    .Z(_02235_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09921_ (.I(_02226_),
    .Z(_02236_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09922_ (.A1(\channels.sus_rel2[4] ),
    .A2(_02236_),
    .B(_02232_),
    .ZN(_02237_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09923_ (.A1(_02234_),
    .A2(_02235_),
    .B(_02237_),
    .ZN(_00217_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09924_ (.I(_02154_),
    .Z(_02238_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09925_ (.A1(\channels.sus_rel2[5] ),
    .A2(_02236_),
    .B(_02232_),
    .ZN(_02239_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09926_ (.A1(_02238_),
    .A2(_02235_),
    .B(_02239_),
    .ZN(_00218_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09927_ (.I(_01813_),
    .Z(_02240_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09928_ (.A1(\channels.sus_rel2[6] ),
    .A2(_02236_),
    .B(_02232_),
    .ZN(_02241_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09929_ (.A1(_02240_),
    .A2(_02235_),
    .B(_02241_),
    .ZN(_00219_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09930_ (.I(_01818_),
    .Z(_02242_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09931_ (.I(_02216_),
    .Z(_02243_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09932_ (.A1(\channels.sus_rel2[7] ),
    .A2(_02236_),
    .B(_02243_),
    .ZN(_02244_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09933_ (.A1(_02242_),
    .A2(_02235_),
    .B(_02244_),
    .ZN(_00220_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09934_ (.I(_02104_),
    .Z(_02245_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09935_ (.A1(_02208_),
    .A2(_01833_),
    .Z(_02246_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09936_ (.I(_02246_),
    .Z(_02247_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09937_ (.I(_02246_),
    .Z(_02248_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09938_ (.A1(\channels.freq3[8] ),
    .A2(_02248_),
    .B(_02243_),
    .ZN(_02249_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09939_ (.A1(_02245_),
    .A2(_02247_),
    .B(_02249_),
    .ZN(_00221_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09940_ (.I(_02184_),
    .Z(_02250_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09941_ (.A1(\channels.freq3[9] ),
    .A2(_02248_),
    .B(_02243_),
    .ZN(_02251_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09942_ (.A1(_02250_),
    .A2(_02247_),
    .B(_02251_),
    .ZN(_00222_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09943_ (.I(_02187_),
    .Z(_02252_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09944_ (.A1(\channels.freq3[10] ),
    .A2(_02248_),
    .B(_02243_),
    .ZN(_02253_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09945_ (.A1(_02252_),
    .A2(_02247_),
    .B(_02253_),
    .ZN(_00223_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09946_ (.I(_02174_),
    .Z(_02254_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09947_ (.I(_02254_),
    .Z(_02255_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09948_ (.A1(\channels.freq3[11] ),
    .A2(_02248_),
    .B(_02255_),
    .ZN(_02256_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09949_ (.A1(_02215_),
    .A2(_02247_),
    .B(_02256_),
    .ZN(_00224_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09950_ (.I(_02246_),
    .Z(_02257_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09951_ (.I(_02246_),
    .Z(_02258_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09952_ (.A1(\channels.freq3[12] ),
    .A2(_02258_),
    .B(_02255_),
    .ZN(_02259_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09953_ (.A1(_02234_),
    .A2(_02257_),
    .B(_02259_),
    .ZN(_00225_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09954_ (.A1(\channels.freq3[13] ),
    .A2(_02258_),
    .B(_02255_),
    .ZN(_02260_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09955_ (.A1(_02238_),
    .A2(_02257_),
    .B(_02260_),
    .ZN(_00226_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09956_ (.A1(\channels.freq3[14] ),
    .A2(_02258_),
    .B(_02255_),
    .ZN(_02261_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09957_ (.A1(_02240_),
    .A2(_02257_),
    .B(_02261_),
    .ZN(_00227_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09958_ (.I(_02254_),
    .Z(_02262_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09959_ (.A1(\channels.freq3[15] ),
    .A2(_02258_),
    .B(_02262_),
    .ZN(_02263_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09960_ (.A1(_02242_),
    .A2(_02257_),
    .B(_02263_),
    .ZN(_00228_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09961_ (.A1(_01781_),
    .A2(_01842_),
    .Z(_02264_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09962_ (.I(_02264_),
    .Z(_02265_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09963_ (.I(_02264_),
    .Z(_02266_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09964_ (.A1(\channels.pw3[8] ),
    .A2(_02266_),
    .B(_02262_),
    .ZN(_02267_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09965_ (.A1(_02245_),
    .A2(_02265_),
    .B(_02267_),
    .ZN(_00229_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09966_ (.A1(\channels.pw3[9] ),
    .A2(_02266_),
    .B(_02262_),
    .ZN(_02268_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09967_ (.A1(_02250_),
    .A2(_02265_),
    .B(_02268_),
    .ZN(_00230_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09968_ (.A1(\channels.pw3[10] ),
    .A2(_02266_),
    .B(_02262_),
    .ZN(_02269_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09969_ (.A1(_02252_),
    .A2(_02265_),
    .B(_02269_),
    .ZN(_00231_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09970_ (.I(\channels.pw3[11] ),
    .ZN(_02270_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09971_ (.A1(_02098_),
    .A2(_02266_),
    .ZN(_02271_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _09972_ (.I(_02101_),
    .Z(_02272_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09973_ (.I(_02272_),
    .Z(_02273_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09974_ (.A1(_02270_),
    .A2(_02265_),
    .B(_02271_),
    .C(_02273_),
    .ZN(_00232_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09975_ (.A1(_02208_),
    .A2(_01881_),
    .Z(_02274_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09976_ (.I(_02274_),
    .Z(_02275_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09977_ (.I(_02274_),
    .Z(_02276_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09978_ (.I(_02254_),
    .Z(_02277_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09979_ (.A1(\channels.ctrl_reg3[0] ),
    .A2(_02276_),
    .B(_02277_),
    .ZN(_02278_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09980_ (.A1(_02245_),
    .A2(_02275_),
    .B(_02278_),
    .ZN(_00233_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09981_ (.A1(\channels.ctrl_reg3[1] ),
    .A2(_02276_),
    .B(_02277_),
    .ZN(_02279_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09982_ (.A1(_02250_),
    .A2(_02275_),
    .B(_02279_),
    .ZN(_00234_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09983_ (.A1(\channels.ctrl_reg3[2] ),
    .A2(_02276_),
    .B(_02277_),
    .ZN(_02280_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09984_ (.A1(_02252_),
    .A2(_02275_),
    .B(_02280_),
    .ZN(_00235_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09985_ (.A1(\channels.ctrl_reg3[3] ),
    .A2(_02276_),
    .B(_02277_),
    .ZN(_02281_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09986_ (.A1(_02215_),
    .A2(_02275_),
    .B(_02281_),
    .ZN(_00236_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09987_ (.I(_02274_),
    .Z(_02282_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09988_ (.I(_02274_),
    .Z(_02283_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09989_ (.I(_02254_),
    .Z(_02284_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09990_ (.A1(\channels.ctrl_reg3[4] ),
    .A2(_02283_),
    .B(_02284_),
    .ZN(_02285_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09991_ (.A1(_02234_),
    .A2(_02282_),
    .B(_02285_),
    .ZN(_00237_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09992_ (.A1(\channels.ctrl_reg3[5] ),
    .A2(_02283_),
    .B(_02284_),
    .ZN(_02286_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09993_ (.A1(_02238_),
    .A2(_02282_),
    .B(_02286_),
    .ZN(_00238_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09994_ (.A1(\channels.ctrl_reg3[6] ),
    .A2(_02283_),
    .B(_02284_),
    .ZN(_02287_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09995_ (.A1(_02240_),
    .A2(_02282_),
    .B(_02287_),
    .ZN(_00239_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09996_ (.A1(\channels.ctrl_reg3[7] ),
    .A2(_02283_),
    .B(_02284_),
    .ZN(_02288_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09997_ (.A1(_02242_),
    .A2(_02282_),
    .B(_02288_),
    .ZN(_00240_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09998_ (.I(_01779_),
    .Z(_02289_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09999_ (.A1(_02289_),
    .A2(_01867_),
    .Z(_02290_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10000_ (.I(_02290_),
    .Z(_02291_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10001_ (.I(_02290_),
    .Z(_02292_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10002_ (.I(_02174_),
    .Z(_02293_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10003_ (.I(_02293_),
    .Z(_02294_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10004_ (.A1(\channels.atk_dec3[0] ),
    .A2(_02292_),
    .B(_02294_),
    .ZN(_02295_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10005_ (.A1(_02245_),
    .A2(_02291_),
    .B(_02295_),
    .ZN(_00241_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10006_ (.A1(\channels.atk_dec3[1] ),
    .A2(_02292_),
    .B(_02294_),
    .ZN(_02296_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10007_ (.A1(_02250_),
    .A2(_02291_),
    .B(_02296_),
    .ZN(_00242_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10008_ (.A1(\channels.atk_dec3[2] ),
    .A2(_02292_),
    .B(_02294_),
    .ZN(_02297_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10009_ (.A1(_02252_),
    .A2(_02291_),
    .B(_02297_),
    .ZN(_00243_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10010_ (.I(_01775_),
    .Z(_02298_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10011_ (.I(_02298_),
    .Z(_02299_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10012_ (.A1(\channels.atk_dec3[3] ),
    .A2(_02292_),
    .B(_02294_),
    .ZN(_02300_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10013_ (.A1(_02299_),
    .A2(_02291_),
    .B(_02300_),
    .ZN(_00244_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10014_ (.I(_02290_),
    .Z(_02301_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10015_ (.I(_02290_),
    .Z(_02302_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10016_ (.I(_02293_),
    .Z(_02303_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10017_ (.A1(\channels.atk_dec3[4] ),
    .A2(_02302_),
    .B(_02303_),
    .ZN(_02304_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10018_ (.A1(_02234_),
    .A2(_02301_),
    .B(_02304_),
    .ZN(_00245_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10019_ (.A1(\channels.atk_dec3[5] ),
    .A2(_02302_),
    .B(_02303_),
    .ZN(_02305_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10020_ (.A1(_02238_),
    .A2(_02301_),
    .B(_02305_),
    .ZN(_00246_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10021_ (.A1(\channels.atk_dec3[6] ),
    .A2(_02302_),
    .B(_02303_),
    .ZN(_02306_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10022_ (.A1(_02240_),
    .A2(_02301_),
    .B(_02306_),
    .ZN(_00247_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10023_ (.A1(\channels.atk_dec3[7] ),
    .A2(_02302_),
    .B(_02303_),
    .ZN(_02307_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10024_ (.A1(_02242_),
    .A2(_02301_),
    .B(_02307_),
    .ZN(_00248_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10025_ (.I(_02104_),
    .Z(_02308_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10026_ (.A1(_02289_),
    .A2(_01943_),
    .Z(_02309_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10027_ (.I(_02309_),
    .Z(_02310_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10028_ (.I(_02309_),
    .Z(_02311_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10029_ (.I(_02293_),
    .Z(_02312_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10030_ (.A1(\channels.sus_rel3[0] ),
    .A2(_02311_),
    .B(_02312_),
    .ZN(_02313_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10031_ (.A1(_02308_),
    .A2(_02310_),
    .B(_02313_),
    .ZN(_00249_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10032_ (.I(_02184_),
    .Z(_02314_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10033_ (.A1(\channels.sus_rel3[1] ),
    .A2(_02311_),
    .B(_02312_),
    .ZN(_02315_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10034_ (.A1(_02314_),
    .A2(_02310_),
    .B(_02315_),
    .ZN(_00250_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10035_ (.I(_02187_),
    .Z(_02316_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10036_ (.A1(\channels.sus_rel3[2] ),
    .A2(_02311_),
    .B(_02312_),
    .ZN(_02317_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10037_ (.A1(_02316_),
    .A2(_02310_),
    .B(_02317_),
    .ZN(_00251_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10038_ (.A1(\channels.sus_rel3[3] ),
    .A2(_02311_),
    .B(_02312_),
    .ZN(_02318_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10039_ (.A1(_02299_),
    .A2(_02310_),
    .B(_02318_),
    .ZN(_00252_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10040_ (.I(_02149_),
    .Z(_02319_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10041_ (.I(_02309_),
    .Z(_02320_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10042_ (.I(_02309_),
    .Z(_02321_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10043_ (.I(_02293_),
    .Z(_02322_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10044_ (.A1(\channels.sus_rel3[4] ),
    .A2(_02321_),
    .B(_02322_),
    .ZN(_02323_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10045_ (.A1(_02319_),
    .A2(_02320_),
    .B(_02323_),
    .ZN(_00253_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10046_ (.I(_02154_),
    .Z(_02324_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10047_ (.A1(\channels.sus_rel3[5] ),
    .A2(_02321_),
    .B(_02322_),
    .ZN(_02325_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10048_ (.A1(_02324_),
    .A2(_02320_),
    .B(_02325_),
    .ZN(_00254_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10049_ (.I(_01813_),
    .Z(_02326_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10050_ (.A1(\channels.sus_rel3[6] ),
    .A2(_02321_),
    .B(_02322_),
    .ZN(_02327_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10051_ (.A1(_02326_),
    .A2(_02320_),
    .B(_02327_),
    .ZN(_00255_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10052_ (.I(_01818_),
    .Z(_02328_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10053_ (.A1(\channels.sus_rel3[7] ),
    .A2(_02321_),
    .B(_02322_),
    .ZN(_02329_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10054_ (.A1(_02328_),
    .A2(_02320_),
    .B(_02329_),
    .ZN(_00256_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10055_ (.A1(_02289_),
    .A2(_01956_),
    .Z(_02330_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10056_ (.I(_02330_),
    .Z(_02331_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10057_ (.I(_02330_),
    .Z(_02332_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10058_ (.I(_01750_),
    .Z(_02333_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10059_ (.I(_02333_),
    .Z(_02334_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10060_ (.I(_02334_),
    .Z(_02335_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10061_ (.A1(\filters.cutoff_lut[9] ),
    .A2(_02332_),
    .B(_02335_),
    .ZN(_02336_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10062_ (.A1(_02308_),
    .A2(_02331_),
    .B(_02336_),
    .ZN(_00257_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10063_ (.A1(\filters.cutoff_lut[10] ),
    .A2(_02332_),
    .B(_02335_),
    .ZN(_02337_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10064_ (.A1(_02314_),
    .A2(_02331_),
    .B(_02337_),
    .ZN(_00258_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10065_ (.A1(\filters.cutoff_lut[11] ),
    .A2(_02332_),
    .B(_02335_),
    .ZN(_02338_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10066_ (.A1(_02316_),
    .A2(_02331_),
    .B(_02338_),
    .ZN(_00259_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10067_ (.A1(\filters.cutoff_lut[12] ),
    .A2(_02332_),
    .B(_02335_),
    .ZN(_02339_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10068_ (.A1(_02299_),
    .A2(_02331_),
    .B(_02339_),
    .ZN(_00260_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10069_ (.I(_02330_),
    .Z(_02340_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10070_ (.I(_02330_),
    .Z(_02341_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10071_ (.I(_02334_),
    .Z(_02342_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10072_ (.A1(\filters.cutoff_lut[13] ),
    .A2(_02341_),
    .B(_02342_),
    .ZN(_02343_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10073_ (.A1(_02319_),
    .A2(_02340_),
    .B(_02343_),
    .ZN(_00261_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10074_ (.A1(\filters.cutoff_lut[14] ),
    .A2(_02341_),
    .B(_02342_),
    .ZN(_02344_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10075_ (.A1(_02324_),
    .A2(_02340_),
    .B(_02344_),
    .ZN(_00262_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10076_ (.A1(\filters.cutoff_lut[15] ),
    .A2(_02341_),
    .B(_02342_),
    .ZN(_02345_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10077_ (.A1(_02326_),
    .A2(_02340_),
    .B(_02345_),
    .ZN(_00263_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10078_ (.A1(\filters.cutoff_lut[16] ),
    .A2(_02341_),
    .B(_02342_),
    .ZN(_02346_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10079_ (.A1(_02328_),
    .A2(_02340_),
    .B(_02346_),
    .ZN(_00264_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10080_ (.I(\tt_um_rejunity_sn76489.chan[2].attenuation.in ),
    .Z(_02347_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _10081_ (.I0(\tt_um_rejunity_sn76489.noise[0].gen.counter[4] ),
    .I1(\tt_um_rejunity_sn76489.noise[0].gen.counter[5] ),
    .I2(\tt_um_rejunity_sn76489.noise[0].gen.counter[6] ),
    .I3(_02347_),
    .S0(\tt_um_rejunity_sn76489.control_noise[0][0] ),
    .S1(\tt_um_rejunity_sn76489.control_noise[0][1] ),
    .Z(_02348_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10082_ (.I(_02348_),
    .ZN(_02349_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10083_ (.A1(_01933_),
    .A2(_02349_),
    .ZN(_00265_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10084_ (.I(\clk_trg[0] ),
    .ZN(_02350_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _10085_ (.A1(_02088_),
    .A2(_01905_),
    .ZN(_02351_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10086_ (.A1(net8),
    .A2(_02351_),
    .ZN(_02352_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10087_ (.I(_01724_),
    .Z(_02353_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10088_ (.I(_02353_),
    .Z(_02354_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _10089_ (.A1(_02350_),
    .A2(_02351_),
    .B(_02352_),
    .C(_02354_),
    .ZN(_00266_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10090_ (.A1(net9),
    .A2(_02351_),
    .ZN(_02355_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _10091_ (.A1(_01065_),
    .A2(_02351_),
    .B(_02355_),
    .C(_02354_),
    .ZN(_00267_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10092_ (.I(_01082_),
    .Z(_02356_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10093_ (.A1(_01070_),
    .A2(_02356_),
    .ZN(_02357_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10094_ (.I(_02357_),
    .Z(_02358_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10095_ (.I(_02358_),
    .Z(_02359_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _10096_ (.I(_01085_),
    .ZN(_02360_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10097_ (.A1(_02360_),
    .A2(_01569_),
    .ZN(_02361_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10098_ (.A1(\channels.sync_outs[2] ),
    .A2(_01245_),
    .ZN(_02362_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10099_ (.A1(_02359_),
    .A2(_02361_),
    .B(_02362_),
    .ZN(_00268_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10100_ (.I(_01282_),
    .Z(_02363_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10101_ (.A1(_01070_),
    .A2(_02363_),
    .ZN(_02364_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10102_ (.I(_02364_),
    .Z(_02365_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10103_ (.I(_02365_),
    .Z(_02366_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10104_ (.A1(\channels.sync_outs[1] ),
    .A2(_01230_),
    .ZN(_02367_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10105_ (.A1(_02366_),
    .A2(_02361_),
    .B(_02367_),
    .ZN(_00269_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10106_ (.A1(\channels.sync_outs[0] ),
    .A2(_01560_),
    .ZN(_02368_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10107_ (.A1(_01540_),
    .A2(_02361_),
    .B(_02368_),
    .ZN(_00270_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10108_ (.A1(_01267_),
    .A2(\channels.ctrl_reg2[4] ),
    .ZN(_02369_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _10109_ (.A1(_01266_),
    .A2(\channels.ctrl_reg3[4] ),
    .B1(\channels.ctrl_reg1[4] ),
    .B2(_01252_),
    .ZN(_02370_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _10110_ (.A1(_01264_),
    .A2(_02369_),
    .B(_02370_),
    .ZN(_02371_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10111_ (.I(_02371_),
    .Z(_02372_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10112_ (.A1(\channels.ctrl_reg2[2] ),
    .A2(\channels.ring_outs[0] ),
    .A3(_01273_),
    .ZN(_02373_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10113_ (.A1(\channels.ctrl_reg3[2] ),
    .A2(\channels.ring_outs[1] ),
    .A3(_01073_),
    .ZN(_02374_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10114_ (.A1(\channels.ctrl_reg1[2] ),
    .A2(\channels.ring_outs[2] ),
    .A3(_01284_),
    .ZN(_02375_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10115_ (.A1(_02373_),
    .A2(_02374_),
    .A3(_02375_),
    .ZN(_02376_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _10116_ (.A1(_02360_),
    .A2(_02376_),
    .Z(_02377_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10117_ (.I(_02377_),
    .Z(_02378_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10118_ (.A1(_01527_),
    .A2(_02378_),
    .Z(_02379_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10119_ (.A1(\channels.ctrl_reg1[5] ),
    .A2(_01286_),
    .Z(_02380_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _10120_ (.A1(\channels.ctrl_reg3[5] ),
    .A2(_01074_),
    .B1(_01274_),
    .B2(\channels.ctrl_reg2[5] ),
    .C(_02380_),
    .ZN(_02381_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10121_ (.I(_02381_),
    .Z(_02382_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10122_ (.A1(\channels.ctrl_reg3[7] ),
    .A2(_01073_),
    .ZN(_02383_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _10123_ (.A1(\channels.ctrl_reg2[7] ),
    .A2(_01273_),
    .B1(_01286_),
    .B2(\channels.ctrl_reg1[7] ),
    .ZN(_02384_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _10124_ (.A1(_02383_),
    .A2(_02384_),
    .ZN(_02385_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10125_ (.I(_02385_),
    .Z(_02386_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10126_ (.A1(_01632_),
    .A2(_02386_),
    .ZN(_02387_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10127_ (.A1(_01534_),
    .A2(_02382_),
    .B(_02387_),
    .ZN(_02388_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10128_ (.I(_01248_),
    .Z(_02389_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10129_ (.I(_01272_),
    .Z(_02390_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10130_ (.A1(_02389_),
    .A2(_02390_),
    .A3(\channels.pw3[11] ),
    .ZN(_02391_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10131_ (.A1(_02390_),
    .A2(\channels.pw2[11] ),
    .B(_01096_),
    .ZN(_02392_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _10132_ (.A1(\channels.pw1[11] ),
    .A2(_01251_),
    .ZN(_02393_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10133_ (.A1(_02391_),
    .A2(_02392_),
    .B(_02393_),
    .ZN(_02394_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _10134_ (.A1(_02360_),
    .A2(_02394_),
    .ZN(_02395_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10135_ (.A1(_02391_),
    .A2(_02392_),
    .Z(_02396_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10136_ (.I(_01071_),
    .Z(_02397_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10137_ (.A1(_02397_),
    .A2(_01250_),
    .A3(\channels.pw2[10] ),
    .ZN(_02398_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10138_ (.A1(_02389_),
    .A2(_02390_),
    .A3(\channels.pw3[10] ),
    .ZN(_02399_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10139_ (.A1(\channels.pw1[10] ),
    .A2(_01285_),
    .ZN(_02400_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _10140_ (.A1(_02398_),
    .A2(_02399_),
    .A3(_02400_),
    .Z(_02401_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _10141_ (.I0(\channels.accum[0][22] ),
    .I1(\channels.accum[1][22] ),
    .I2(\channels.accum[2][22] ),
    .I3(\channels.accum[3][22] ),
    .S0(_01495_),
    .S1(_01496_),
    .Z(_02402_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _10142_ (.A1(_01085_),
    .A2(_02396_),
    .A3(_02393_),
    .B1(_02401_),
    .B2(_02402_),
    .ZN(_02403_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10143_ (.I(_01555_),
    .ZN(_02404_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10144_ (.I(_01272_),
    .Z(_02405_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10145_ (.A1(_02389_),
    .A2(_02405_),
    .A3(\channels.pw3[9] ),
    .ZN(_02406_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10146_ (.A1(_02390_),
    .A2(\channels.pw2[9] ),
    .B(_02397_),
    .ZN(_02407_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10147_ (.A1(\channels.pw1[9] ),
    .A2(_01251_),
    .ZN(_02408_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10148_ (.A1(_02406_),
    .A2(_02407_),
    .B(_02408_),
    .ZN(_02409_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10149_ (.A1(_02397_),
    .A2(_01250_),
    .A3(\channels.pw2[8] ),
    .ZN(_02410_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10150_ (.A1(_02389_),
    .A2(_02405_),
    .A3(\channels.pw3[8] ),
    .ZN(_02411_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10151_ (.A1(\channels.pw1[8] ),
    .A2(_01285_),
    .ZN(_02412_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10152_ (.A1(_02410_),
    .A2(_02411_),
    .A3(_02412_),
    .ZN(_02413_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10153_ (.A1(_02404_),
    .A2(_02409_),
    .B1(_02413_),
    .B2(_01553_),
    .ZN(_02414_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10154_ (.A1(_02398_),
    .A2(_02399_),
    .A3(_02400_),
    .ZN(_02415_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _10155_ (.A1(_01566_),
    .A2(_02415_),
    .B1(_02409_),
    .B2(_02404_),
    .ZN(_02416_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10156_ (.A1(_02414_),
    .A2(_02416_),
    .ZN(_02417_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _10157_ (.A1(_02403_),
    .A2(_02417_),
    .ZN(_02418_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10158_ (.A1(_02406_),
    .A2(_02407_),
    .Z(_02419_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _10159_ (.A1(_02410_),
    .A2(_02411_),
    .A3(_02412_),
    .Z(_02420_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _10160_ (.A1(_01555_),
    .A2(_02419_),
    .A3(_02408_),
    .B1(_02420_),
    .B2(_01550_),
    .ZN(_02421_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10161_ (.A1(_02360_),
    .A2(_02394_),
    .B1(_02413_),
    .B2(_01553_),
    .ZN(_02422_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _10162_ (.A1(_02403_),
    .A2(_02421_),
    .A3(_02416_),
    .A4(_02422_),
    .ZN(_02423_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10163_ (.I(_02423_),
    .ZN(_02424_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _10164_ (.A1(_01097_),
    .A2(_01098_),
    .A3(\channels.pw2[7] ),
    .ZN(_02425_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10165_ (.I(_01249_),
    .Z(_02426_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10166_ (.I(_01272_),
    .Z(_02427_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10167_ (.I(_02427_),
    .Z(_02428_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _10168_ (.A1(_02426_),
    .A2(_02428_),
    .A3(\channels.pw3[7] ),
    .ZN(_02429_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10169_ (.I(_01284_),
    .Z(_02430_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _10170_ (.A1(\channels.pw1[7] ),
    .A2(_02430_),
    .ZN(_02431_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _10171_ (.A1(_01541_),
    .A2(_02425_),
    .A3(_02429_),
    .A4(_02431_),
    .ZN(_02432_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _10172_ (.A1(_02425_),
    .A2(_02429_),
    .A3(_02431_),
    .Z(_02433_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _10173_ (.I(\channels.pw1[5] ),
    .ZN(_02434_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10174_ (.I(_01285_),
    .Z(_02435_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _10175_ (.A1(_02426_),
    .A2(_02405_),
    .A3(\channels.pw3[5] ),
    .ZN(_02436_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10176_ (.A1(_02428_),
    .A2(\channels.pw2[5] ),
    .B(_01097_),
    .ZN(_02437_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _10177_ (.A1(_02434_),
    .A2(_02435_),
    .B1(_02436_),
    .B2(_02437_),
    .C(_01527_),
    .ZN(_02438_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _10178_ (.I(\channels.pw1[4] ),
    .ZN(_02439_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _10179_ (.A1(_02426_),
    .A2(_02428_),
    .A3(\channels.pw3[4] ),
    .ZN(_02440_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10180_ (.A1(_02428_),
    .A2(\channels.pw2[4] ),
    .B(_01097_),
    .ZN(_02441_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _10181_ (.A1(_02439_),
    .A2(_01286_),
    .B1(_02440_),
    .B2(_02441_),
    .C(_01520_),
    .ZN(_02442_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _10182_ (.A1(_02438_),
    .A2(_02442_),
    .ZN(_02443_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _10183_ (.A1(_02397_),
    .A2(_01098_),
    .A3(\channels.pw2[6] ),
    .ZN(_02444_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _10184_ (.A1(_02426_),
    .A2(_02405_),
    .A3(\channels.pw3[6] ),
    .ZN(_02445_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10185_ (.A1(\channels.pw1[6] ),
    .A2(_02430_),
    .ZN(_02446_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _10186_ (.A1(_01533_),
    .A2(_02444_),
    .A3(_02445_),
    .A4(_02446_),
    .ZN(_02447_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10187_ (.A1(_01265_),
    .A2(_01263_),
    .A3(\channels.pw2[5] ),
    .ZN(_02448_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10188_ (.A1(\channels.pw1[5] ),
    .A2(_02435_),
    .ZN(_02449_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _10189_ (.A1(_01527_),
    .A2(_02448_),
    .A3(_02436_),
    .A4(_02449_),
    .ZN(_02450_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _10190_ (.A1(_02447_),
    .A2(_02450_),
    .ZN(_02451_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _10191_ (.A1(_02444_),
    .A2(_02445_),
    .A3(_02446_),
    .Z(_02452_));
 gf180mcu_fd_sc_mcu7t5v0__oai222_4 _10192_ (.A1(_01541_),
    .A2(_02433_),
    .B1(_02443_),
    .B2(_02451_),
    .C1(_02452_),
    .C2(_01533_),
    .ZN(_02453_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10193_ (.I(\channels.pw2[2] ),
    .ZN(_02454_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10194_ (.I(_02427_),
    .Z(_02455_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10195_ (.A1(_01582_),
    .A2(_02455_),
    .A3(\channels.pw3[2] ),
    .ZN(_02456_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10196_ (.A1(\channels.pw1[2] ),
    .A2(_02430_),
    .ZN(_02457_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _10197_ (.A1(_02454_),
    .A2(_01099_),
    .B(_02456_),
    .C(_02457_),
    .ZN(_02458_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10198_ (.A1(_01498_),
    .A2(_02458_),
    .ZN(_02459_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _10199_ (.A1(_01265_),
    .A2(_01263_),
    .A3(\channels.pw2[0] ),
    .ZN(_02460_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10200_ (.A1(_01582_),
    .A2(_02455_),
    .A3(\channels.pw3[0] ),
    .ZN(_02461_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10201_ (.A1(\channels.pw1[0] ),
    .A2(_02435_),
    .ZN(_02462_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _10202_ (.A1(_01469_),
    .A2(_02460_),
    .A3(_02461_),
    .A4(_02462_),
    .ZN(_02463_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _10203_ (.A1(_01249_),
    .A2(_02427_),
    .A3(\channels.pw3[1] ),
    .ZN(_02464_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10204_ (.A1(_01072_),
    .A2(\channels.pw1[1] ),
    .Z(_02465_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _10205_ (.A1(_02427_),
    .A2(\channels.pw2[1] ),
    .B(_02465_),
    .C(_01096_),
    .ZN(_02466_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10206_ (.A1(_01481_),
    .A2(_02464_),
    .A3(_02466_),
    .ZN(_02467_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10207_ (.A1(_02464_),
    .A2(_02466_),
    .B(_01481_),
    .ZN(_02468_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10208_ (.A1(_02463_),
    .A2(_02467_),
    .B(_02468_),
    .ZN(_02469_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10209_ (.I(\channels.pw2[3] ),
    .ZN(_02470_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _10210_ (.A1(_01582_),
    .A2(_02455_),
    .A3(\channels.pw3[3] ),
    .ZN(_02471_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10211_ (.A1(\channels.pw1[3] ),
    .A2(_02430_),
    .ZN(_02472_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _10212_ (.A1(_02470_),
    .A2(_01099_),
    .B(_02471_),
    .C(_02472_),
    .ZN(_02473_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10213_ (.A1(_01509_),
    .A2(_02473_),
    .B1(_02458_),
    .B2(_01498_),
    .ZN(_02474_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10214_ (.A1(_02459_),
    .A2(_02469_),
    .B(_02474_),
    .ZN(_02475_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_4 _10215_ (.A1(_01541_),
    .A2(_02433_),
    .B1(_02452_),
    .B2(_01533_),
    .ZN(_02476_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10216_ (.A1(_02438_),
    .A2(_02442_),
    .Z(_02477_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10217_ (.A1(_01265_),
    .A2(_01098_),
    .A3(\channels.pw2[4] ),
    .ZN(_02478_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10218_ (.A1(\channels.pw1[4] ),
    .A2(_02435_),
    .ZN(_02479_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _10219_ (.A1(_01520_),
    .A2(_02478_),
    .A3(_02440_),
    .A4(_02479_),
    .ZN(_02480_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10220_ (.A1(_01509_),
    .A2(_02473_),
    .B(_02480_),
    .C(_02432_),
    .ZN(_02481_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _10221_ (.A1(_02476_),
    .A2(_02477_),
    .A3(_02451_),
    .A4(_02481_),
    .ZN(_02482_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _10222_ (.A1(_02432_),
    .A2(_02453_),
    .B1(_02475_),
    .B2(_02482_),
    .ZN(_02483_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_4 _10223_ (.A1(_02395_),
    .A2(_02418_),
    .B1(_02424_),
    .B2(_02483_),
    .ZN(_02484_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10224_ (.A1(_02432_),
    .A2(_02480_),
    .ZN(_02485_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _10225_ (.A1(_02476_),
    .A2(_02477_),
    .A3(_02451_),
    .A4(_02485_),
    .ZN(_02486_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10226_ (.A1(_02464_),
    .A2(_02466_),
    .ZN(_02487_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10227_ (.A1(_01481_),
    .A2(_02487_),
    .ZN(_02488_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10228_ (.A1(_02463_),
    .A2(_02488_),
    .Z(_02489_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10229_ (.A1(_01510_),
    .A2(_02473_),
    .ZN(_02490_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10230_ (.A1(_02461_),
    .A2(_02462_),
    .Z(_02491_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10231_ (.A1(_02460_),
    .A2(_02491_),
    .B(_01469_),
    .ZN(_02492_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _10232_ (.A1(_02459_),
    .A2(_02490_),
    .A3(_02492_),
    .ZN(_02493_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _10233_ (.A1(_02423_),
    .A2(_02474_),
    .A3(_02489_),
    .A4(_02493_),
    .Z(_02494_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10234_ (.A1(_01266_),
    .A2(\channels.ctrl_reg2[6] ),
    .ZN(_02495_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10235_ (.A1(_01263_),
    .A2(_02495_),
    .ZN(_02496_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _10236_ (.A1(_01266_),
    .A2(\channels.ctrl_reg3[6] ),
    .B1(\channels.ctrl_reg1[6] ),
    .B2(_01252_),
    .C(_02496_),
    .ZN(_02497_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _10237_ (.A1(_02486_),
    .A2(_02494_),
    .B(_02497_),
    .ZN(_02498_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _10238_ (.A1(_02484_),
    .A2(_02498_),
    .Z(_02499_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _10239_ (.A1(_02372_),
    .A2(_02379_),
    .B(_02388_),
    .C(_02499_),
    .ZN(_02500_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10240_ (.I(_02500_),
    .Z(_02501_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10241_ (.I(_02501_),
    .Z(_02502_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _10242_ (.I0(\channels.env_vol[0][0] ),
    .I1(\channels.env_vol[1][0] ),
    .I2(\channels.ch3_env[0] ),
    .I3(\channels.env_vol[3][0] ),
    .S0(_01145_),
    .S1(_01159_),
    .Z(_02503_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10243_ (.I(_02503_),
    .Z(_02504_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10244_ (.I(_02504_),
    .Z(_02505_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10245_ (.A1(_02502_),
    .A2(_02505_),
    .Z(_02506_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10246_ (.A1(_02484_),
    .A2(_02498_),
    .B(_02386_),
    .ZN(_02507_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10247_ (.I(_02507_),
    .Z(_02508_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10248_ (.I(_02508_),
    .Z(_02509_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10249_ (.A1(_01497_),
    .A2(_02378_),
    .Z(_02510_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10250_ (.A1(_01508_),
    .A2(_02381_),
    .ZN(_02511_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10251_ (.A1(_02372_),
    .A2(_02510_),
    .B(_02511_),
    .ZN(_02512_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10252_ (.I(_02512_),
    .Z(_02513_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10253_ (.I(_02513_),
    .Z(_02514_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10254_ (.I(\channels.ch3_env[2] ),
    .ZN(_02515_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10255_ (.A1(_01306_),
    .A2(_02515_),
    .ZN(_02516_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10256_ (.A1(_01306_),
    .A2(\channels.env_vol[3][2] ),
    .B(_02516_),
    .ZN(_02517_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10257_ (.I(_01141_),
    .Z(_02518_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10258_ (.I(_02518_),
    .Z(_02519_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10259_ (.I0(\channels.env_vol[0][2] ),
    .I1(\channels.env_vol[1][2] ),
    .S(_02519_),
    .Z(_02520_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10260_ (.A1(_01157_),
    .A2(_02520_),
    .ZN(_02521_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10261_ (.A1(_01688_),
    .A2(_02517_),
    .B(_02521_),
    .ZN(_02522_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _10262_ (.A1(_02509_),
    .A2(_02514_),
    .A3(_02522_),
    .Z(_02523_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10263_ (.I(_02508_),
    .Z(_02524_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10264_ (.A1(_01482_),
    .A2(_02378_),
    .Z(_02525_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10265_ (.A1(_01497_),
    .A2(_02382_),
    .ZN(_02526_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10266_ (.A1(_02372_),
    .A2(_02525_),
    .B(_02526_),
    .ZN(_02527_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10267_ (.I(_02527_),
    .Z(_02528_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10268_ (.I(_01656_),
    .Z(_02529_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10269_ (.I(\channels.ch3_env[3] ),
    .ZN(_02530_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10270_ (.A1(_01305_),
    .A2(_02530_),
    .ZN(_02531_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10271_ (.A1(_01143_),
    .A2(\channels.env_vol[3][3] ),
    .B(_02531_),
    .ZN(_02532_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10272_ (.I0(\channels.env_vol[0][3] ),
    .I1(\channels.env_vol[1][3] ),
    .S(_02518_),
    .Z(_02533_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10273_ (.A1(_01156_),
    .A2(_02533_),
    .ZN(_02534_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10274_ (.A1(_02529_),
    .A2(_02532_),
    .B(_02534_),
    .ZN(_02535_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10275_ (.I(_02535_),
    .Z(_02536_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _10276_ (.A1(_02524_),
    .A2(_02528_),
    .A3(_02536_),
    .ZN(_02537_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _10277_ (.I(_02372_),
    .Z(_02538_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10278_ (.I(_02378_),
    .Z(_02539_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10279_ (.A1(_01470_),
    .A2(_02539_),
    .Z(_02540_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10280_ (.I(_02382_),
    .Z(_02541_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10281_ (.A1(_01482_),
    .A2(_02541_),
    .ZN(_02542_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _10282_ (.A1(_02538_),
    .A2(_02540_),
    .B(_02542_),
    .ZN(_02543_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _10283_ (.I0(\channels.env_vol[0][4] ),
    .I1(\channels.env_vol[1][4] ),
    .I2(\channels.ch3_env[4] ),
    .I3(\channels.env_vol[3][4] ),
    .S0(_01143_),
    .S1(_01687_),
    .Z(_02544_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _10284_ (.A1(_02524_),
    .A2(_02543_),
    .A3(_02544_),
    .ZN(_02545_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10285_ (.A1(_02537_),
    .A2(_02545_),
    .ZN(_02546_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10286_ (.A1(_02537_),
    .A2(_02545_),
    .ZN(_02547_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10287_ (.A1(_02523_),
    .A2(_02546_),
    .B(_02547_),
    .ZN(_02548_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10288_ (.A1(_01521_),
    .A2(_02377_),
    .ZN(_02549_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10289_ (.I(_02371_),
    .ZN(_02550_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10290_ (.A1(_01615_),
    .A2(_02385_),
    .ZN(_02551_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _10291_ (.A1(_01528_),
    .A2(_02382_),
    .B1(_02549_),
    .B2(_02550_),
    .C(_02551_),
    .ZN(_02552_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10292_ (.A1(_02484_),
    .A2(_02498_),
    .B(_02552_),
    .ZN(_02553_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10293_ (.I(_02553_),
    .Z(_02554_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10294_ (.I(_02554_),
    .Z(_02555_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10295_ (.I(\channels.ch3_env[1] ),
    .ZN(_02556_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10296_ (.A1(_01307_),
    .A2(_02556_),
    .ZN(_02557_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10297_ (.A1(_01307_),
    .A2(\channels.env_vol[3][1] ),
    .B(_02557_),
    .ZN(_02558_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10298_ (.I0(\channels.env_vol[0][1] ),
    .I1(\channels.env_vol[1][1] ),
    .S(_01144_),
    .Z(_02559_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10299_ (.A1(_01328_),
    .A2(_02559_),
    .ZN(_02560_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10300_ (.A1(_01328_),
    .A2(_02558_),
    .B(_02560_),
    .ZN(_02561_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10301_ (.I(_02561_),
    .Z(_02562_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10302_ (.A1(_02555_),
    .A2(_02562_),
    .ZN(_02563_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10303_ (.A1(_02548_),
    .A2(_02563_),
    .ZN(_02564_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10304_ (.A1(_02548_),
    .A2(_02563_),
    .ZN(_02565_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10305_ (.A1(_02506_),
    .A2(_02564_),
    .B(_02565_),
    .ZN(_02566_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10306_ (.I(_02539_),
    .Z(_02567_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10307_ (.A1(_01470_),
    .A2(_02541_),
    .ZN(_02568_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _10308_ (.A1(_02567_),
    .A2(_02538_),
    .B(_02568_),
    .ZN(_02569_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10309_ (.I(\channels.ch3_env[6] ),
    .ZN(_02570_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10310_ (.A1(_02518_),
    .A2(_02570_),
    .ZN(_02571_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10311_ (.A1(_02519_),
    .A2(\channels.env_vol[3][6] ),
    .B(_02571_),
    .ZN(_02572_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10312_ (.I0(\channels.env_vol[0][6] ),
    .I1(\channels.env_vol[1][6] ),
    .S(_01142_),
    .Z(_02573_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10313_ (.A1(_01156_),
    .A2(_02573_),
    .ZN(_02574_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10314_ (.A1(_01687_),
    .A2(_02572_),
    .B(_02574_),
    .ZN(_02575_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10315_ (.I(_02575_),
    .Z(_02576_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _10316_ (.A1(_02524_),
    .A2(_02569_),
    .A3(_02576_),
    .ZN(_02577_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10317_ (.I(\channels.ch3_env[5] ),
    .ZN(_02578_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10318_ (.A1(_01143_),
    .A2(_02578_),
    .ZN(_02579_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10319_ (.A1(_01306_),
    .A2(\channels.env_vol[3][5] ),
    .B(_02579_),
    .ZN(_02580_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10320_ (.I0(\channels.env_vol[0][5] ),
    .I1(\channels.env_vol[1][5] ),
    .S(_02519_),
    .Z(_02581_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10321_ (.A1(_01157_),
    .A2(_02581_),
    .ZN(_02582_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10322_ (.A1(_01688_),
    .A2(_02580_),
    .B(_02582_),
    .ZN(_02583_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _10323_ (.A1(_02524_),
    .A2(_02543_),
    .A3(_02583_),
    .ZN(_02584_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10324_ (.A1(_02577_),
    .A2(_02584_),
    .ZN(_02585_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10325_ (.A1(_01510_),
    .A2(_02377_),
    .Z(_02586_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10326_ (.A1(_01598_),
    .A2(_02385_),
    .ZN(_02587_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _10327_ (.A1(_01521_),
    .A2(_02381_),
    .B1(_02586_),
    .B2(_02550_),
    .C(_02587_),
    .ZN(_02588_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10328_ (.A1(_02484_),
    .A2(_02498_),
    .B(_02588_),
    .ZN(_02589_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10329_ (.I(_02589_),
    .Z(_02590_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10330_ (.A1(_02522_),
    .A2(_02590_),
    .ZN(_02591_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10331_ (.I(_02507_),
    .Z(_02592_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _10332_ (.A1(_02592_),
    .A2(_02535_),
    .A3(_02513_),
    .ZN(_02593_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10333_ (.I(_02544_),
    .Z(_02594_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _10334_ (.A1(_02509_),
    .A2(_02528_),
    .A3(_02594_),
    .ZN(_02595_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _10335_ (.A1(_02591_),
    .A2(_02593_),
    .A3(_02595_),
    .Z(_02596_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10336_ (.A1(_02585_),
    .A2(_02596_),
    .Z(_02597_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10337_ (.I(_02592_),
    .Z(_02598_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10338_ (.I(_02598_),
    .Z(_02599_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10339_ (.I(_02569_),
    .Z(_02600_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10340_ (.I(_02583_),
    .Z(_02601_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10341_ (.I(_02601_),
    .Z(_02602_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _10342_ (.A1(_02599_),
    .A2(_02600_),
    .A3(_02602_),
    .ZN(_02603_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _10343_ (.A1(_02537_),
    .A2(_02545_),
    .A3(_02523_),
    .ZN(_02604_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10344_ (.A1(_02603_),
    .A2(_02604_),
    .ZN(_02605_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10345_ (.A1(_02597_),
    .A2(_02605_),
    .ZN(_02606_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10346_ (.I(_02503_),
    .Z(_02607_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10347_ (.A1(_02502_),
    .A2(_02607_),
    .ZN(_02608_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _10348_ (.A1(_02548_),
    .A2(_02563_),
    .A3(_02608_),
    .Z(_02609_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10349_ (.A1(_02597_),
    .A2(_02605_),
    .ZN(_02610_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10350_ (.A1(_02606_),
    .A2(_02609_),
    .B(_02610_),
    .ZN(_02611_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10351_ (.A1(_02585_),
    .A2(_02596_),
    .ZN(_02612_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10352_ (.I(_02591_),
    .ZN(_02613_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10353_ (.A1(_02593_),
    .A2(_02595_),
    .ZN(_02614_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10354_ (.A1(_02593_),
    .A2(_02595_),
    .ZN(_02615_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10355_ (.A1(_02613_),
    .A2(_02614_),
    .B(_02615_),
    .ZN(_02616_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10356_ (.A1(_02562_),
    .A2(_02502_),
    .ZN(_02617_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10357_ (.A1(_02616_),
    .A2(_02617_),
    .Z(_02618_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10358_ (.A1(_01534_),
    .A2(_02539_),
    .Z(_02619_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10359_ (.A1(_01657_),
    .A2(_02386_),
    .ZN(_02620_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10360_ (.A1(_01542_),
    .A2(_02541_),
    .B(_02620_),
    .ZN(_02621_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _10361_ (.A1(_02538_),
    .A2(_02619_),
    .B(_02621_),
    .C(_02499_),
    .ZN(_02622_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10362_ (.I(_02622_),
    .Z(_02623_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10363_ (.I(_02623_),
    .Z(_02624_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10364_ (.A1(_02504_),
    .A2(_02624_),
    .ZN(_02625_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10365_ (.A1(_02618_),
    .A2(_02625_),
    .Z(_02626_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10366_ (.A1(_02577_),
    .A2(_02584_),
    .ZN(_02627_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10367_ (.I(_02528_),
    .Z(_02628_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10368_ (.A1(_02598_),
    .A2(_02628_),
    .A3(_02601_),
    .ZN(_02629_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10369_ (.I(_02543_),
    .Z(_02630_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _10370_ (.A1(_02598_),
    .A2(_02630_),
    .A3(_02576_),
    .ZN(_02631_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10371_ (.I(\channels.ch3_env[7] ),
    .ZN(_02632_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10372_ (.A1(_01305_),
    .A2(_02632_),
    .ZN(_02633_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10373_ (.A1(_02519_),
    .A2(\channels.env_vol[3][7] ),
    .B(_02633_),
    .ZN(_02634_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10374_ (.I0(\channels.env_vol[0][7] ),
    .I1(\channels.env_vol[1][7] ),
    .S(_02518_),
    .Z(_02635_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10375_ (.A1(_01156_),
    .A2(_02635_),
    .ZN(_02636_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10376_ (.A1(_02529_),
    .A2(_02634_),
    .B(_02636_),
    .ZN(_02637_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10377_ (.I(_02637_),
    .Z(_02638_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _10378_ (.A1(_02509_),
    .A2(_02569_),
    .A3(_02638_),
    .ZN(_02639_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _10379_ (.A1(_02629_),
    .A2(_02631_),
    .A3(_02639_),
    .ZN(_02640_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10380_ (.I(_02522_),
    .Z(_02641_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10381_ (.I(_02641_),
    .Z(_02642_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10382_ (.A1(_02642_),
    .A2(_02555_),
    .ZN(_02643_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10383_ (.I(_02536_),
    .Z(_02644_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10384_ (.I(_02590_),
    .Z(_02645_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10385_ (.A1(_02644_),
    .A2(_02645_),
    .ZN(_02646_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10386_ (.A1(_02509_),
    .A2(_02594_),
    .A3(_02513_),
    .ZN(_02647_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10387_ (.A1(_02646_),
    .A2(_02647_),
    .ZN(_02648_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10388_ (.A1(_02643_),
    .A2(_02648_),
    .ZN(_02649_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _10389_ (.A1(_02627_),
    .A2(_02640_),
    .A3(_02649_),
    .ZN(_02650_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _10390_ (.A1(_02612_),
    .A2(_02626_),
    .A3(_02650_),
    .ZN(_02651_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _10391_ (.A1(_02566_),
    .A2(_02611_),
    .A3(_02651_),
    .ZN(_02652_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10392_ (.A1(_02555_),
    .A2(_02503_),
    .Z(_02653_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _10393_ (.A1(_02599_),
    .A2(_02628_),
    .A3(_02642_),
    .ZN(_02654_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10394_ (.I(_02598_),
    .Z(_02655_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _10395_ (.A1(_02655_),
    .A2(_02644_),
    .A3(_02630_),
    .ZN(_02656_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10396_ (.I(_02544_),
    .Z(_02657_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _10397_ (.A1(_02655_),
    .A2(_02657_),
    .A3(_02569_),
    .ZN(_02658_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10398_ (.A1(_02656_),
    .A2(_02658_),
    .Z(_02659_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10399_ (.A1(_02656_),
    .A2(_02658_),
    .Z(_02660_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10400_ (.A1(_02654_),
    .A2(_02659_),
    .B(_02660_),
    .ZN(_02661_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10401_ (.I(_02561_),
    .Z(_02662_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10402_ (.A1(_02662_),
    .A2(_02645_),
    .Z(_02663_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10403_ (.A1(_02661_),
    .A2(_02663_),
    .Z(_02664_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10404_ (.A1(_02661_),
    .A2(_02663_),
    .Z(_02665_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10405_ (.A1(_02653_),
    .A2(_02664_),
    .B(_02665_),
    .ZN(_02666_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10406_ (.A1(_02603_),
    .A2(_02604_),
    .Z(_02667_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _10407_ (.A1(_02653_),
    .A2(_02661_),
    .A3(_02663_),
    .Z(_02668_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10408_ (.A1(_02667_),
    .A2(_02668_),
    .Z(_02669_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10409_ (.A1(_02606_),
    .A2(_02609_),
    .Z(_02670_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10410_ (.A1(_02669_),
    .A2(_02670_),
    .ZN(_02671_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10411_ (.A1(_02669_),
    .A2(_02670_),
    .ZN(_02672_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10412_ (.A1(_02666_),
    .A2(_02671_),
    .B(_02672_),
    .ZN(_02673_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10413_ (.A1(_02667_),
    .A2(_02668_),
    .ZN(_02674_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10414_ (.A1(_02599_),
    .A2(_02514_),
    .A3(_02662_),
    .ZN(_02675_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10415_ (.I(_02644_),
    .Z(_02676_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _10416_ (.A1(_02655_),
    .A2(_02676_),
    .A3(_02600_),
    .ZN(_02677_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _10417_ (.A1(_02655_),
    .A2(_02630_),
    .A3(_02641_),
    .ZN(_02678_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _10418_ (.A1(_02677_),
    .A2(_02678_),
    .ZN(_02679_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10419_ (.A1(_02607_),
    .A2(_02645_),
    .ZN(_02680_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _10420_ (.A1(_02675_),
    .A2(_02679_),
    .A3(_02680_),
    .ZN(_02681_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _10421_ (.A1(_02656_),
    .A2(_02658_),
    .A3(_02654_),
    .Z(_02682_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _10422_ (.A1(_02669_),
    .A2(_02674_),
    .A3(_02681_),
    .A4(_02682_),
    .ZN(_02683_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10423_ (.I(_02599_),
    .Z(_02684_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10424_ (.I(_02684_),
    .Z(_02685_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10425_ (.I(_02562_),
    .Z(_02686_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10426_ (.I(_02686_),
    .Z(_02687_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _10427_ (.A1(_02685_),
    .A2(_02514_),
    .A3(_02687_),
    .A4(_02679_),
    .ZN(_02688_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10428_ (.A1(_02675_),
    .A2(_02679_),
    .Z(_02689_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10429_ (.A1(_02689_),
    .A2(_02680_),
    .Z(_02690_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10430_ (.A1(_02681_),
    .A2(_02682_),
    .ZN(_02691_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _10431_ (.A1(_02667_),
    .A2(_02668_),
    .A3(_02691_),
    .ZN(_02692_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10432_ (.A1(_02688_),
    .A2(_02690_),
    .B(_02692_),
    .ZN(_02693_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _10433_ (.A1(_02669_),
    .A2(_02670_),
    .A3(_02666_),
    .ZN(_02694_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10434_ (.A1(_02683_),
    .A2(_02693_),
    .B(_02694_),
    .ZN(_02695_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10435_ (.A1(_02681_),
    .A2(_02682_),
    .Z(_02696_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10436_ (.A1(_02684_),
    .A2(_02628_),
    .A3(_02686_),
    .ZN(_02697_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10437_ (.A1(_02684_),
    .A2(_02514_),
    .A3(_02607_),
    .ZN(_02698_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10438_ (.A1(_02697_),
    .A2(_02698_),
    .ZN(_02699_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10439_ (.A1(_02677_),
    .A2(_02678_),
    .ZN(_02700_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10440_ (.A1(_02697_),
    .A2(_02698_),
    .Z(_02701_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10441_ (.A1(_02699_),
    .A2(_02700_),
    .B(_02701_),
    .ZN(_02702_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10442_ (.I(_02505_),
    .Z(_02703_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10443_ (.A1(_02684_),
    .A2(_02630_),
    .ZN(_02704_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10444_ (.A1(_01162_),
    .A2(_02558_),
    .ZN(_02705_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10445_ (.A1(_01162_),
    .A2(_02559_),
    .B(_02705_),
    .ZN(_02706_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10446_ (.I(_02706_),
    .Z(_02707_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10447_ (.A1(_02704_),
    .A2(_02707_),
    .ZN(_02708_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _10448_ (.A1(_02685_),
    .A2(_02628_),
    .A3(_02703_),
    .A4(_02708_),
    .ZN(_02709_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10449_ (.I(_02642_),
    .Z(_02710_));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 _10450_ (.I(_02505_),
    .ZN(_02711_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10451_ (.A1(_02508_),
    .A2(_02527_),
    .ZN(_02712_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10452_ (.I(_02712_),
    .Z(_02713_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10453_ (.A1(_02704_),
    .A2(_02706_),
    .B1(_02711_),
    .B2(_02713_),
    .ZN(_02714_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _10454_ (.A1(_02685_),
    .A2(_02710_),
    .A3(_02600_),
    .A4(_02714_),
    .ZN(_02715_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10455_ (.A1(_02699_),
    .A2(_02700_),
    .ZN(_02716_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10456_ (.A1(_02709_),
    .A2(_02715_),
    .B(_02716_),
    .ZN(_02717_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _10457_ (.A1(_02681_),
    .A2(_02682_),
    .A3(_02702_),
    .Z(_02718_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10458_ (.A1(_02717_),
    .A2(_02718_),
    .Z(_02719_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10459_ (.A1(_01164_),
    .A2(_02517_),
    .ZN(_02720_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10460_ (.A1(_01164_),
    .A2(_02520_),
    .B(_02720_),
    .ZN(_02721_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10461_ (.A1(_02713_),
    .A2(_02721_),
    .B(_02716_),
    .ZN(_02722_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _10462_ (.A1(_02685_),
    .A2(_02703_),
    .A3(_02600_),
    .A4(_02708_),
    .ZN(_02723_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10463_ (.A1(_02654_),
    .A2(_02716_),
    .Z(_02724_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10464_ (.A1(_02717_),
    .A2(_02718_),
    .ZN(_02725_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _10465_ (.A1(_02722_),
    .A2(_02723_),
    .A3(_02724_),
    .B(_02725_),
    .ZN(_02726_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10466_ (.A1(_02696_),
    .A2(_02702_),
    .B1(_02719_),
    .B2(_02726_),
    .ZN(_02727_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10467_ (.A1(_02688_),
    .A2(_02690_),
    .A3(_02692_),
    .ZN(_02728_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _10468_ (.A1(_02683_),
    .A2(_02693_),
    .A3(_02694_),
    .B(_02728_),
    .ZN(_02729_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _10469_ (.A1(_02693_),
    .A2(_02727_),
    .A3(_02729_),
    .Z(_02730_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10470_ (.A1(_02652_),
    .A2(_02673_),
    .ZN(_02731_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10471_ (.A1(_02695_),
    .A2(_02730_),
    .B(_02731_),
    .ZN(_02732_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10472_ (.A1(_02652_),
    .A2(_02673_),
    .B(_02732_),
    .ZN(_02733_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10473_ (.A1(_02611_),
    .A2(_02651_),
    .ZN(_02734_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10474_ (.A1(_02611_),
    .A2(_02651_),
    .ZN(_02735_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10475_ (.A1(_02566_),
    .A2(_02734_),
    .B(_02735_),
    .ZN(_02736_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10476_ (.A1(_02703_),
    .A2(_02618_),
    .A3(_02624_),
    .ZN(_02737_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10477_ (.A1(_02616_),
    .A2(_02617_),
    .B(_02737_),
    .ZN(_02738_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10478_ (.A1(_02612_),
    .A2(_02650_),
    .ZN(_02739_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10479_ (.A1(_02612_),
    .A2(_02650_),
    .ZN(_02740_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10480_ (.A1(_02626_),
    .A2(_02739_),
    .B(_02740_),
    .ZN(_02741_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10481_ (.A1(_02627_),
    .A2(_02640_),
    .ZN(_02742_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10482_ (.A1(_02627_),
    .A2(_02640_),
    .ZN(_02743_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10483_ (.A1(_02742_),
    .A2(_02649_),
    .B(_02743_),
    .ZN(_02744_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10484_ (.A1(_02631_),
    .A2(_02639_),
    .Z(_02745_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10485_ (.A1(_02631_),
    .A2(_02639_),
    .Z(_02746_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10486_ (.A1(_02629_),
    .A2(_02745_),
    .B(_02746_),
    .ZN(_02747_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _10487_ (.A1(_02592_),
    .A2(_02543_),
    .A3(_02638_),
    .ZN(_02748_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _10488_ (.A1(_02592_),
    .A2(_02528_),
    .A3(_02576_),
    .ZN(_02749_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10489_ (.A1(_02507_),
    .A2(_02512_),
    .ZN(_02750_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10490_ (.A1(_01688_),
    .A2(_02580_),
    .ZN(_02751_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _10491_ (.A1(_01158_),
    .A2(_02581_),
    .B(_02751_),
    .ZN(_02752_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10492_ (.A1(_02750_),
    .A2(_02752_),
    .ZN(_02753_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _10493_ (.A1(_02748_),
    .A2(_02749_),
    .A3(_02753_),
    .Z(_02754_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10494_ (.A1(_02641_),
    .A2(_02501_),
    .ZN(_02755_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10495_ (.A1(_02594_),
    .A2(_02645_),
    .ZN(_02756_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10496_ (.A1(_02536_),
    .A2(_02554_),
    .ZN(_02757_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10497_ (.A1(_02756_),
    .A2(_02757_),
    .Z(_02758_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10498_ (.A1(_02756_),
    .A2(_02757_),
    .ZN(_02759_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10499_ (.A1(_02758_),
    .A2(_02759_),
    .ZN(_02760_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10500_ (.A1(_02755_),
    .A2(_02760_),
    .Z(_02761_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _10501_ (.A1(_02747_),
    .A2(_02754_),
    .A3(_02761_),
    .Z(_02762_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10502_ (.A1(_02744_),
    .A2(_02762_),
    .ZN(_02763_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10503_ (.A1(_02646_),
    .A2(_02647_),
    .Z(_02764_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10504_ (.A1(_02643_),
    .A2(_02648_),
    .B(_02764_),
    .ZN(_02765_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10505_ (.A1(_02662_),
    .A2(_02623_),
    .ZN(_02766_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10506_ (.A1(_02765_),
    .A2(_02766_),
    .Z(_02767_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _10507_ (.I(_02538_),
    .Z(_02768_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10508_ (.A1(_01542_),
    .A2(_02539_),
    .Z(_02769_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10509_ (.I(_02541_),
    .Z(_02770_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10510_ (.I(_02386_),
    .Z(_02771_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10511_ (.A1(_01668_),
    .A2(_02771_),
    .ZN(_02772_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10512_ (.A1(_01550_),
    .A2(_02770_),
    .B(_02772_),
    .ZN(_02773_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _10513_ (.I(_02499_),
    .Z(_02774_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _10514_ (.A1(_02768_),
    .A2(_02769_),
    .B(_02773_),
    .C(_02774_),
    .ZN(_02775_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10515_ (.I(_02775_),
    .Z(_02776_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10516_ (.I(_02776_),
    .Z(_02777_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10517_ (.A1(_02504_),
    .A2(_02777_),
    .ZN(_02778_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10518_ (.A1(_02767_),
    .A2(_02778_),
    .ZN(_02779_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10519_ (.A1(_02763_),
    .A2(_02779_),
    .Z(_02780_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10520_ (.A1(_02741_),
    .A2(_02780_),
    .Z(_02781_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10521_ (.A1(_02738_),
    .A2(_02781_),
    .Z(_02782_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _10522_ (.A1(_02733_),
    .A2(_02736_),
    .A3(_02782_),
    .Z(_02783_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10523_ (.I(_01089_),
    .Z(_02784_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10524_ (.A1(\channels.sample3[0] ),
    .A2(_02784_),
    .ZN(_02785_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10525_ (.A1(_02359_),
    .A2(_02783_),
    .B(_02785_),
    .ZN(_00271_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10526_ (.A1(_02736_),
    .A2(_02782_),
    .ZN(_02786_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10527_ (.A1(_02736_),
    .A2(_02782_),
    .ZN(_02787_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10528_ (.A1(_02733_),
    .A2(_02786_),
    .B(_02787_),
    .ZN(_02788_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10529_ (.A1(_02741_),
    .A2(_02780_),
    .Z(_02789_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10530_ (.A1(_02738_),
    .A2(_02781_),
    .B(_02789_),
    .ZN(_02790_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10531_ (.A1(_02686_),
    .A2(_02624_),
    .A3(_02765_),
    .ZN(_02791_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10532_ (.A1(_02767_),
    .A2(_02778_),
    .B(_02791_),
    .ZN(_02792_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10533_ (.A1(_02744_),
    .A2(_02762_),
    .ZN(_02793_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10534_ (.A1(_02763_),
    .A2(_02779_),
    .B(_02793_),
    .ZN(_02794_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10535_ (.A1(_02747_),
    .A2(_02754_),
    .Z(_02795_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10536_ (.A1(_02747_),
    .A2(_02754_),
    .Z(_02796_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10537_ (.A1(_02795_),
    .A2(_02761_),
    .B(_02796_),
    .ZN(_02797_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10538_ (.A1(_02748_),
    .A2(_02749_),
    .ZN(_02798_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10539_ (.A1(_02748_),
    .A2(_02749_),
    .ZN(_02799_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10540_ (.A1(_02798_),
    .A2(_02753_),
    .B(_02799_),
    .ZN(_02800_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10541_ (.A1(_02529_),
    .A2(_02634_),
    .ZN(_02801_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10542_ (.A1(_01157_),
    .A2(_02635_),
    .B(_02801_),
    .ZN(_02802_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10543_ (.A1(_02712_),
    .A2(_02802_),
    .ZN(_02803_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10544_ (.A1(_01687_),
    .A2(_02572_),
    .ZN(_02804_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10545_ (.A1(_02529_),
    .A2(_02573_),
    .B(_02804_),
    .ZN(_02805_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10546_ (.A1(_02750_),
    .A2(_02805_),
    .ZN(_02806_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10547_ (.A1(_02583_),
    .A2(_02590_),
    .Z(_02807_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _10548_ (.A1(_02803_),
    .A2(_02806_),
    .A3(_02807_),
    .ZN(_02808_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10549_ (.A1(_02800_),
    .A2(_02808_),
    .Z(_02809_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10550_ (.A1(_02522_),
    .A2(_02622_),
    .ZN(_02810_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10551_ (.A1(_02544_),
    .A2(_02554_),
    .ZN(_02811_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10552_ (.A1(_02535_),
    .A2(_02500_),
    .ZN(_02812_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10553_ (.A1(_02811_),
    .A2(_02812_),
    .ZN(_02813_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10554_ (.A1(_02810_),
    .A2(_02813_),
    .Z(_02814_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10555_ (.A1(_02809_),
    .A2(_02814_),
    .ZN(_02815_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10556_ (.A1(_02797_),
    .A2(_02815_),
    .Z(_02816_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10557_ (.A1(_02755_),
    .A2(_02760_),
    .B(_02758_),
    .ZN(_02817_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10558_ (.A1(_02561_),
    .A2(_02776_),
    .ZN(_02818_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10559_ (.A1(_02817_),
    .A2(_02818_),
    .ZN(_02819_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10560_ (.A1(_01550_),
    .A2(_02567_),
    .Z(_02820_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10561_ (.A1(_01689_),
    .A2(_02771_),
    .ZN(_02821_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10562_ (.A1(_01556_),
    .A2(_02770_),
    .B(_02821_),
    .ZN(_02822_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _10563_ (.A1(_02768_),
    .A2(_02820_),
    .B(_02822_),
    .C(_02774_),
    .ZN(_02823_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10564_ (.I(_02823_),
    .Z(_02824_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10565_ (.A1(_02607_),
    .A2(_02824_),
    .ZN(_02825_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10566_ (.A1(_02819_),
    .A2(_02825_),
    .ZN(_02826_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10567_ (.A1(_02816_),
    .A2(_02826_),
    .Z(_02827_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10568_ (.A1(_02794_),
    .A2(_02827_),
    .Z(_02828_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10569_ (.A1(_02792_),
    .A2(_02828_),
    .ZN(_02829_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10570_ (.A1(_02790_),
    .A2(_02829_),
    .ZN(_02830_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _10571_ (.A1(_02788_),
    .A2(_02830_),
    .Z(_02831_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10572_ (.A1(\channels.sample3[1] ),
    .A2(_02784_),
    .ZN(_02832_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10573_ (.A1(_02359_),
    .A2(_02831_),
    .B(_02832_),
    .ZN(_00272_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10574_ (.I(_02830_),
    .ZN(_02833_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10575_ (.A1(_02790_),
    .A2(_02829_),
    .ZN(_02834_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10576_ (.A1(_02788_),
    .A2(_02833_),
    .B(_02834_),
    .ZN(_02835_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10577_ (.A1(_02794_),
    .A2(_02827_),
    .Z(_02836_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10578_ (.A1(_02792_),
    .A2(_02828_),
    .B(_02836_),
    .ZN(_02837_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10579_ (.A1(_02687_),
    .A2(_02777_),
    .A3(_02817_),
    .ZN(_02838_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10580_ (.I(_02703_),
    .Z(_02839_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10581_ (.I(_02824_),
    .Z(_02840_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10582_ (.A1(_02839_),
    .A2(_02819_),
    .A3(_02840_),
    .ZN(_02841_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10583_ (.A1(_02838_),
    .A2(_02841_),
    .Z(_02842_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10584_ (.A1(_02797_),
    .A2(_02815_),
    .ZN(_02843_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10585_ (.A1(_02816_),
    .A2(_02826_),
    .B(_02843_),
    .ZN(_02844_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10586_ (.A1(_02800_),
    .A2(_02808_),
    .ZN(_02845_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10587_ (.A1(_02809_),
    .A2(_02814_),
    .B(_02845_),
    .ZN(_02846_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10588_ (.I(_02802_),
    .Z(_02847_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10589_ (.A1(_02750_),
    .A2(_02805_),
    .B1(_02847_),
    .B2(_02713_),
    .ZN(_02848_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _10590_ (.A1(_02713_),
    .A2(_02750_),
    .A3(_02805_),
    .A4(_02847_),
    .ZN(_02849_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10591_ (.A1(_02848_),
    .A2(_02807_),
    .B(_02849_),
    .ZN(_02850_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10592_ (.A1(_02554_),
    .A2(_02601_),
    .ZN(_02851_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10593_ (.A1(_02508_),
    .A2(_02513_),
    .A3(_02637_),
    .ZN(_02852_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10594_ (.A1(_02575_),
    .A2(_02589_),
    .ZN(_02853_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10595_ (.A1(_02852_),
    .A2(_02853_),
    .ZN(_02854_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10596_ (.A1(_02851_),
    .A2(_02854_),
    .ZN(_02855_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10597_ (.A1(_02850_),
    .A2(_02855_),
    .Z(_02856_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10598_ (.A1(_02850_),
    .A2(_02855_),
    .ZN(_02857_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10599_ (.A1(_02856_),
    .A2(_02857_),
    .ZN(_02858_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10600_ (.A1(_02641_),
    .A2(_02775_),
    .ZN(_02859_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10601_ (.A1(_02594_),
    .A2(_02500_),
    .ZN(_02860_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10602_ (.A1(_02536_),
    .A2(_02622_),
    .ZN(_02861_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10603_ (.A1(_02860_),
    .A2(_02861_),
    .ZN(_02862_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10604_ (.A1(_02859_),
    .A2(_02862_),
    .ZN(_02863_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10605_ (.A1(_02858_),
    .A2(_02863_),
    .ZN(_02864_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10606_ (.A1(_02811_),
    .A2(_02812_),
    .Z(_02865_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10607_ (.A1(_02810_),
    .A2(_02813_),
    .B(_02865_),
    .ZN(_02866_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10608_ (.A1(_02562_),
    .A2(_02823_),
    .ZN(_02867_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10609_ (.A1(_02866_),
    .A2(_02867_),
    .ZN(_02868_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10610_ (.A1(_01556_),
    .A2(_02567_),
    .Z(_02869_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10611_ (.A1(_01705_),
    .A2(_02771_),
    .ZN(_02870_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10612_ (.A1(_02402_),
    .A2(_02770_),
    .B(_02870_),
    .ZN(_02871_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _10613_ (.A1(_02768_),
    .A2(_02869_),
    .B(_02871_),
    .C(_02774_),
    .ZN(_02872_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10614_ (.I(_02872_),
    .Z(_02873_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10615_ (.A1(_02504_),
    .A2(_02873_),
    .ZN(_02874_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10616_ (.A1(_02868_),
    .A2(_02874_),
    .ZN(_02875_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _10617_ (.A1(_02846_),
    .A2(_02864_),
    .A3(_02875_),
    .ZN(_02876_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10618_ (.A1(_02844_),
    .A2(_02876_),
    .ZN(_02877_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10619_ (.A1(_02842_),
    .A2(_02877_),
    .ZN(_02878_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10620_ (.A1(_02837_),
    .A2(_02878_),
    .Z(_02879_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _10621_ (.A1(_02835_),
    .A2(_02879_),
    .Z(_02880_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10622_ (.A1(\channels.sample3[2] ),
    .A2(_02784_),
    .ZN(_02881_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10623_ (.A1(_02359_),
    .A2(_02880_),
    .B(_02881_),
    .ZN(_00273_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10624_ (.I(_02358_),
    .Z(_02882_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10625_ (.I(_02879_),
    .ZN(_02883_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10626_ (.A1(_02837_),
    .A2(_02878_),
    .Z(_02884_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10627_ (.A1(_02835_),
    .A2(_02883_),
    .B(_02884_),
    .ZN(_02885_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10628_ (.A1(_02844_),
    .A2(_02876_),
    .ZN(_02886_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10629_ (.A1(_02842_),
    .A2(_02877_),
    .ZN(_02887_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10630_ (.A1(_02886_),
    .A2(_02887_),
    .ZN(_02888_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10631_ (.A1(_02687_),
    .A2(_02840_),
    .A3(_02866_),
    .ZN(_02889_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10632_ (.I(_02873_),
    .Z(_02890_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10633_ (.A1(_02839_),
    .A2(_02868_),
    .A3(_02890_),
    .ZN(_02891_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10634_ (.A1(_02889_),
    .A2(_02891_),
    .Z(_02892_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10635_ (.A1(_02846_),
    .A2(_02864_),
    .ZN(_02893_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10636_ (.A1(_02846_),
    .A2(_02864_),
    .ZN(_02894_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10637_ (.A1(_02893_),
    .A2(_02875_),
    .B(_02894_),
    .ZN(_02895_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10638_ (.A1(_02858_),
    .A2(_02863_),
    .B(_02856_),
    .ZN(_02896_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10639_ (.A1(_02852_),
    .A2(_02853_),
    .ZN(_02897_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10640_ (.A1(_02851_),
    .A2(_02854_),
    .ZN(_02898_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10641_ (.A1(_02897_),
    .A2(_02898_),
    .ZN(_02899_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10642_ (.A1(_02501_),
    .A2(_02601_),
    .ZN(_02900_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10643_ (.A1(_02590_),
    .A2(_02637_),
    .ZN(_02901_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10644_ (.A1(_02553_),
    .A2(_02575_),
    .ZN(_02902_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10645_ (.A1(_02901_),
    .A2(_02902_),
    .ZN(_02903_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10646_ (.A1(_02900_),
    .A2(_02903_),
    .Z(_02904_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10647_ (.A1(_02900_),
    .A2(_02903_),
    .ZN(_02905_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10648_ (.A1(_02904_),
    .A2(_02905_),
    .ZN(_02906_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10649_ (.A1(_02899_),
    .A2(_02906_),
    .ZN(_02907_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10650_ (.A1(_02642_),
    .A2(_02823_),
    .ZN(_02908_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10651_ (.A1(_02657_),
    .A2(_02622_),
    .ZN(_02909_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10652_ (.A1(_02644_),
    .A2(_02775_),
    .ZN(_02910_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10653_ (.A1(_02909_),
    .A2(_02910_),
    .ZN(_02911_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10654_ (.A1(_02908_),
    .A2(_02911_),
    .ZN(_02912_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10655_ (.A1(_02907_),
    .A2(_02912_),
    .Z(_02913_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10656_ (.A1(_02896_),
    .A2(_02913_),
    .Z(_02914_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10657_ (.A1(_02860_),
    .A2(_02861_),
    .ZN(_02915_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10658_ (.A1(_02859_),
    .A2(_02862_),
    .ZN(_02916_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10659_ (.A1(_02915_),
    .A2(_02916_),
    .ZN(_02917_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10660_ (.A1(_02662_),
    .A2(_02872_),
    .ZN(_02918_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10661_ (.A1(_02917_),
    .A2(_02918_),
    .Z(_02919_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10662_ (.A1(_02402_),
    .A2(_02567_),
    .Z(_02920_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10663_ (.A1(_01715_),
    .A2(_02771_),
    .ZN(_02921_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10664_ (.A1(_01085_),
    .A2(_02770_),
    .B(_02921_),
    .ZN(_02922_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _10665_ (.A1(_02768_),
    .A2(_02920_),
    .B(_02922_),
    .C(_02774_),
    .ZN(_02923_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10666_ (.A1(_02505_),
    .A2(_02923_),
    .ZN(_02924_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10667_ (.A1(_02919_),
    .A2(_02924_),
    .ZN(_02925_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10668_ (.A1(_02914_),
    .A2(_02925_),
    .ZN(_02926_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10669_ (.A1(_02895_),
    .A2(_02926_),
    .ZN(_02927_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10670_ (.A1(_02892_),
    .A2(_02927_),
    .Z(_02928_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10671_ (.A1(_02892_),
    .A2(_02927_),
    .ZN(_02929_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10672_ (.A1(_02928_),
    .A2(_02929_),
    .ZN(_02930_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10673_ (.A1(_02888_),
    .A2(_02930_),
    .ZN(_02931_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _10674_ (.A1(_02885_),
    .A2(_02931_),
    .Z(_02932_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10675_ (.A1(\channels.sample3[3] ),
    .A2(_02784_),
    .ZN(_02933_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10676_ (.A1(_02882_),
    .A2(_02932_),
    .B(_02933_),
    .ZN(_00274_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10677_ (.I(_02931_),
    .ZN(_02934_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10678_ (.A1(_02888_),
    .A2(_02930_),
    .ZN(_02935_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10679_ (.A1(_02885_),
    .A2(_02934_),
    .B(_02935_),
    .ZN(_02936_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10680_ (.A1(_02895_),
    .A2(_02926_),
    .B(_02928_),
    .ZN(_02937_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10681_ (.A1(_02917_),
    .A2(_02918_),
    .Z(_02938_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10682_ (.I(_02923_),
    .Z(_02939_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10683_ (.I(_02939_),
    .Z(_02940_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10684_ (.A1(_02839_),
    .A2(_02919_),
    .A3(_02940_),
    .ZN(_02941_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10685_ (.A1(_02938_),
    .A2(_02941_),
    .Z(_02942_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10686_ (.A1(_02896_),
    .A2(_02913_),
    .Z(_02943_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10687_ (.A1(_02914_),
    .A2(_02925_),
    .B(_02943_),
    .ZN(_02944_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10688_ (.A1(_02909_),
    .A2(_02910_),
    .ZN(_02945_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10689_ (.A1(_02908_),
    .A2(_02911_),
    .ZN(_02946_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10690_ (.A1(_02945_),
    .A2(_02946_),
    .ZN(_02947_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10691_ (.A1(_02686_),
    .A2(_02923_),
    .ZN(_02948_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10692_ (.A1(_02947_),
    .A2(_02948_),
    .Z(_02949_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10693_ (.A1(_02899_),
    .A2(_02906_),
    .Z(_02950_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10694_ (.A1(_02907_),
    .A2(_02912_),
    .B(_02950_),
    .ZN(_02951_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10695_ (.A1(_02901_),
    .A2(_02902_),
    .B(_02904_),
    .ZN(_02952_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10696_ (.A1(_02602_),
    .A2(_02623_),
    .ZN(_02953_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10697_ (.A1(_02555_),
    .A2(_02638_),
    .ZN(_02954_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10698_ (.I(_02576_),
    .Z(_02955_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10699_ (.A1(_02501_),
    .A2(_02955_),
    .ZN(_02956_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10700_ (.A1(_02954_),
    .A2(_02956_),
    .ZN(_02957_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10701_ (.A1(_02953_),
    .A2(_02957_),
    .Z(_02958_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10702_ (.A1(_02952_),
    .A2(_02958_),
    .Z(_02959_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10703_ (.A1(_02710_),
    .A2(_02873_),
    .ZN(_02960_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10704_ (.I(_02657_),
    .Z(_02961_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10705_ (.A1(_02961_),
    .A2(_02777_),
    .ZN(_02962_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10706_ (.A1(_02676_),
    .A2(_02824_),
    .ZN(_02963_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10707_ (.A1(_02962_),
    .A2(_02963_),
    .Z(_02964_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10708_ (.A1(_02962_),
    .A2(_02963_),
    .ZN(_02965_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10709_ (.A1(_02964_),
    .A2(_02965_),
    .ZN(_02966_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10710_ (.A1(_02960_),
    .A2(_02966_),
    .Z(_02967_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10711_ (.A1(_02959_),
    .A2(_02967_),
    .Z(_02968_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _10712_ (.A1(_02949_),
    .A2(_02951_),
    .A3(_02968_),
    .ZN(_02969_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10713_ (.A1(_02944_),
    .A2(_02969_),
    .ZN(_02970_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10714_ (.A1(_02942_),
    .A2(_02970_),
    .Z(_02971_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10715_ (.A1(_02937_),
    .A2(_02971_),
    .Z(_02972_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _10716_ (.A1(_02936_),
    .A2(_02972_),
    .Z(_02973_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10717_ (.I(_01088_),
    .Z(_02974_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10718_ (.I(_02974_),
    .Z(_02975_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10719_ (.A1(\channels.sample3[4] ),
    .A2(_02975_),
    .ZN(_02976_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10720_ (.A1(_02882_),
    .A2(_02973_),
    .B(_02976_),
    .ZN(_00275_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10721_ (.I(_02972_),
    .ZN(_02977_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10722_ (.A1(_02937_),
    .A2(_02971_),
    .ZN(_02978_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10723_ (.A1(_02936_),
    .A2(_02977_),
    .B(_02978_),
    .ZN(_02979_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10724_ (.A1(_02944_),
    .A2(_02969_),
    .ZN(_02980_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10725_ (.A1(_02942_),
    .A2(_02970_),
    .ZN(_02981_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10726_ (.A1(_02980_),
    .A2(_02981_),
    .ZN(_02982_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10727_ (.A1(_02947_),
    .A2(_02948_),
    .Z(_02983_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10728_ (.A1(_02951_),
    .A2(_02968_),
    .Z(_02984_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10729_ (.A1(_02951_),
    .A2(_02968_),
    .Z(_02985_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10730_ (.A1(_02949_),
    .A2(_02984_),
    .B(_02985_),
    .ZN(_02986_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10731_ (.A1(_02960_),
    .A2(_02966_),
    .B(_02964_),
    .ZN(_02987_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10732_ (.A1(_02952_),
    .A2(_02958_),
    .ZN(_02988_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10733_ (.A1(_02959_),
    .A2(_02967_),
    .ZN(_02989_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10734_ (.A1(_02988_),
    .A2(_02989_),
    .ZN(_02990_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10735_ (.A1(_02953_),
    .A2(_02957_),
    .Z(_02991_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10736_ (.A1(_02954_),
    .A2(_02956_),
    .B(_02991_),
    .ZN(_02992_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10737_ (.A1(_02602_),
    .A2(_02776_),
    .ZN(_02993_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10738_ (.I(_02638_),
    .Z(_02994_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10739_ (.A1(_02502_),
    .A2(_02994_),
    .ZN(_02995_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10740_ (.A1(_02955_),
    .A2(_02623_),
    .ZN(_02996_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10741_ (.A1(_02995_),
    .A2(_02996_),
    .ZN(_02997_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10742_ (.A1(_02993_),
    .A2(_02997_),
    .Z(_02998_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10743_ (.A1(_02992_),
    .A2(_02998_),
    .Z(_02999_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10744_ (.A1(_02710_),
    .A2(_02923_),
    .ZN(_03000_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10745_ (.A1(_02657_),
    .A2(_02823_),
    .ZN(_03001_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10746_ (.A1(_02676_),
    .A2(_02872_),
    .ZN(_03002_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10747_ (.A1(_03001_),
    .A2(_03002_),
    .ZN(_03003_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10748_ (.A1(_03000_),
    .A2(_03003_),
    .Z(_03004_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10749_ (.A1(_02999_),
    .A2(_03004_),
    .Z(_03005_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10750_ (.A1(_02990_),
    .A2(_03005_),
    .Z(_03006_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10751_ (.A1(_02987_),
    .A2(_03006_),
    .ZN(_03007_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10752_ (.A1(_02986_),
    .A2(_03007_),
    .Z(_03008_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10753_ (.A1(_02986_),
    .A2(_03007_),
    .ZN(_03009_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10754_ (.A1(_03008_),
    .A2(_03009_),
    .ZN(_03010_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10755_ (.A1(_02983_),
    .A2(_03010_),
    .Z(_03011_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10756_ (.A1(_02982_),
    .A2(_03011_),
    .Z(_03012_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _10757_ (.A1(_02979_),
    .A2(_03012_),
    .Z(_03013_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10758_ (.A1(_01927_),
    .A2(_02975_),
    .ZN(_03014_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10759_ (.A1(_02882_),
    .A2(_03013_),
    .B(_03014_),
    .ZN(_00276_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10760_ (.A1(_02980_),
    .A2(_02981_),
    .B(_03011_),
    .ZN(_03015_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10761_ (.I(_03012_),
    .ZN(_03016_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10762_ (.A1(_02979_),
    .A2(_03016_),
    .ZN(_03017_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10763_ (.A1(_03015_),
    .A2(_03017_),
    .ZN(_03018_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10764_ (.A1(_02990_),
    .A2(_03005_),
    .ZN(_03019_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10765_ (.A1(_02987_),
    .A2(_03006_),
    .ZN(_03020_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10766_ (.A1(_03001_),
    .A2(_03002_),
    .ZN(_03021_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10767_ (.A1(_03000_),
    .A2(_03003_),
    .ZN(_03022_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10768_ (.A1(_02992_),
    .A2(_02998_),
    .ZN(_03023_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10769_ (.A1(_02999_),
    .A2(_03004_),
    .ZN(_03024_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10770_ (.A1(_03023_),
    .A2(_03024_),
    .ZN(_03025_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10771_ (.A1(_02993_),
    .A2(_02997_),
    .Z(_03026_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10772_ (.A1(_02995_),
    .A2(_02996_),
    .B(_03026_),
    .ZN(_03027_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10773_ (.I(_02602_),
    .Z(_03028_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10774_ (.A1(_03028_),
    .A2(_02840_),
    .ZN(_03029_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10775_ (.A1(_02624_),
    .A2(_02994_),
    .ZN(_03030_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10776_ (.I(_02955_),
    .Z(_03031_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10777_ (.A1(_03031_),
    .A2(_02777_),
    .ZN(_03032_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10778_ (.A1(_03030_),
    .A2(_03032_),
    .Z(_03033_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10779_ (.A1(_03030_),
    .A2(_03032_),
    .ZN(_03034_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10780_ (.A1(_03033_),
    .A2(_03034_),
    .ZN(_03035_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10781_ (.A1(_03029_),
    .A2(_03035_),
    .Z(_03036_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10782_ (.A1(_03027_),
    .A2(_03036_),
    .Z(_03037_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10783_ (.A1(_02961_),
    .A2(_02873_),
    .ZN(_03038_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10784_ (.I(_02676_),
    .Z(_03039_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10785_ (.A1(_03039_),
    .A2(_02939_),
    .ZN(_03040_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10786_ (.A1(_03038_),
    .A2(_03040_),
    .Z(_03041_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10787_ (.A1(_03037_),
    .A2(_03041_),
    .Z(_03042_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10788_ (.A1(_03025_),
    .A2(_03042_),
    .Z(_03043_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10789_ (.A1(_03021_),
    .A2(_03022_),
    .B(_03043_),
    .ZN(_03044_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _10790_ (.A1(_03021_),
    .A2(_03022_),
    .A3(_03043_),
    .Z(_03045_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10791_ (.A1(_03044_),
    .A2(_03045_),
    .ZN(_03046_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10792_ (.A1(_03019_),
    .A2(_03020_),
    .B(_03046_),
    .ZN(_03047_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _10793_ (.A1(_03019_),
    .A2(_03020_),
    .A3(_03046_),
    .Z(_03048_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10794_ (.A1(_03047_),
    .A2(_03048_),
    .ZN(_03049_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10795_ (.A1(_02983_),
    .A2(_03010_),
    .B(_03008_),
    .ZN(_03050_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10796_ (.A1(_03049_),
    .A2(_03050_),
    .ZN(_03051_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _10797_ (.A1(_03018_),
    .A2(_03051_),
    .Z(_03052_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10798_ (.A1(\channels.sample3[6] ),
    .A2(_02975_),
    .ZN(_03053_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10799_ (.A1(_02882_),
    .A2(_03052_),
    .B(_03053_),
    .ZN(_00277_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10800_ (.I(_02358_),
    .Z(_03054_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10801_ (.A1(_03049_),
    .A2(_03050_),
    .Z(_03055_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10802_ (.A1(_03015_),
    .A2(_03017_),
    .B(_03051_),
    .ZN(_03056_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10803_ (.A1(_03055_),
    .A2(_03056_),
    .ZN(_03057_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10804_ (.A1(_03038_),
    .A2(_03040_),
    .Z(_03058_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10805_ (.A1(_03027_),
    .A2(_03036_),
    .ZN(_03059_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10806_ (.A1(_03037_),
    .A2(_03041_),
    .ZN(_03060_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10807_ (.A1(_03059_),
    .A2(_03060_),
    .ZN(_03061_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10808_ (.A1(_02961_),
    .A2(_02939_),
    .ZN(_03062_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10809_ (.A1(_03029_),
    .A2(_03035_),
    .B(_03033_),
    .ZN(_03063_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10810_ (.A1(_03028_),
    .A2(_02872_),
    .ZN(_03064_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10811_ (.A1(_02994_),
    .A2(_02776_),
    .ZN(_03065_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10812_ (.A1(_02955_),
    .A2(_02824_),
    .ZN(_03066_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10813_ (.A1(_03065_),
    .A2(_03066_),
    .Z(_03067_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10814_ (.A1(_03065_),
    .A2(_03066_),
    .ZN(_03068_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10815_ (.A1(_03067_),
    .A2(_03068_),
    .ZN(_03069_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10816_ (.A1(_03064_),
    .A2(_03069_),
    .Z(_03070_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10817_ (.A1(_03063_),
    .A2(_03070_),
    .Z(_03071_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10818_ (.A1(_03062_),
    .A2(_03071_),
    .ZN(_03072_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10819_ (.A1(_03061_),
    .A2(_03072_),
    .ZN(_03073_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10820_ (.A1(_03058_),
    .A2(_03073_),
    .ZN(_03074_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10821_ (.A1(_03025_),
    .A2(_03042_),
    .ZN(_03075_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10822_ (.A1(_03075_),
    .A2(_03044_),
    .Z(_03076_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10823_ (.A1(_03074_),
    .A2(_03076_),
    .ZN(_03077_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10824_ (.A1(_03047_),
    .A2(_03077_),
    .Z(_03078_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10825_ (.I(_03078_),
    .ZN(_03079_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _10826_ (.A1(_03057_),
    .A2(_03079_),
    .Z(_03080_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10827_ (.A1(_01977_),
    .A2(_02975_),
    .ZN(_03081_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10828_ (.A1(_03054_),
    .A2(_03080_),
    .B(_03081_),
    .ZN(_00278_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10829_ (.I(_03077_),
    .ZN(_03082_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10830_ (.A1(_03047_),
    .A2(_03082_),
    .ZN(_03083_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10831_ (.A1(_03055_),
    .A2(_03056_),
    .B(_03079_),
    .ZN(_03084_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10832_ (.A1(_03083_),
    .A2(_03084_),
    .Z(_03085_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10833_ (.A1(_03074_),
    .A2(_03076_),
    .ZN(_03086_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10834_ (.A1(_03028_),
    .A2(_02939_),
    .ZN(_03087_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10835_ (.I(_02994_),
    .Z(_03088_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10836_ (.A1(_03088_),
    .A2(_02840_),
    .ZN(_03089_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10837_ (.A1(_03031_),
    .A2(_02890_),
    .ZN(_03090_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _10838_ (.A1(_03087_),
    .A2(_03089_),
    .A3(_03090_),
    .Z(_03091_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10839_ (.A1(_03064_),
    .A2(_03069_),
    .B(_03067_),
    .ZN(_03092_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10840_ (.I(_03092_),
    .ZN(_03093_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10841_ (.A1(_03091_),
    .A2(_03093_),
    .Z(_03094_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10842_ (.A1(_03063_),
    .A2(_03070_),
    .ZN(_03095_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10843_ (.I(_02961_),
    .Z(_03096_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10844_ (.A1(_03096_),
    .A2(_02940_),
    .A3(_03071_),
    .ZN(_03097_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10845_ (.A1(_03095_),
    .A2(_03097_),
    .ZN(_03098_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10846_ (.A1(_03094_),
    .A2(_03098_),
    .Z(_03099_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10847_ (.A1(_03061_),
    .A2(_03072_),
    .ZN(_03100_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10848_ (.A1(_03058_),
    .A2(_03073_),
    .B(_03100_),
    .ZN(_03101_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10849_ (.A1(_03099_),
    .A2(_03101_),
    .Z(_03102_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10850_ (.A1(_03086_),
    .A2(_03102_),
    .ZN(_03103_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _10851_ (.A1(_03085_),
    .A2(_03103_),
    .ZN(_03104_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10852_ (.I(_02974_),
    .Z(_03105_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10853_ (.A1(\channels.sample3[8] ),
    .A2(_03105_),
    .ZN(_03106_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10854_ (.A1(_03054_),
    .A2(_03104_),
    .B(_03106_),
    .ZN(_00279_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10855_ (.A1(_03086_),
    .A2(_03102_),
    .ZN(_03107_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10856_ (.A1(_03085_),
    .A2(_03103_),
    .B(_03107_),
    .ZN(_03108_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10857_ (.A1(_03099_),
    .A2(_03101_),
    .ZN(_03109_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10858_ (.A1(_03089_),
    .A2(_03090_),
    .Z(_03110_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10859_ (.A1(_03089_),
    .A2(_03090_),
    .Z(_03111_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10860_ (.A1(_03087_),
    .A2(_03110_),
    .B(_03111_),
    .ZN(_03112_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10861_ (.A1(_03088_),
    .A2(_02890_),
    .ZN(_03113_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10862_ (.A1(_03031_),
    .A2(_02940_),
    .ZN(_03114_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10863_ (.A1(_03113_),
    .A2(_03114_),
    .Z(_03115_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10864_ (.A1(_03112_),
    .A2(_03115_),
    .Z(_03116_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10865_ (.A1(_03091_),
    .A2(_03093_),
    .ZN(_03117_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10866_ (.A1(_03094_),
    .A2(_03098_),
    .Z(_03118_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10867_ (.A1(_03117_),
    .A2(_03118_),
    .ZN(_03119_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10868_ (.A1(_03116_),
    .A2(_03119_),
    .Z(_03120_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10869_ (.A1(_03109_),
    .A2(_03120_),
    .Z(_03121_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _10870_ (.A1(_03108_),
    .A2(_03121_),
    .ZN(_03122_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10871_ (.A1(_02029_),
    .A2(_03105_),
    .ZN(_03123_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10872_ (.A1(_03054_),
    .A2(_03122_),
    .B(_03123_),
    .ZN(_00280_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10873_ (.A1(_03108_),
    .A2(_03121_),
    .ZN(_03124_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10874_ (.A1(_03109_),
    .A2(_03120_),
    .B(_03124_),
    .ZN(_03125_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10875_ (.A1(_03118_),
    .A2(_03116_),
    .ZN(_03126_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10876_ (.A1(_03117_),
    .A2(_03116_),
    .ZN(_03127_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10877_ (.I(_03031_),
    .Z(_03128_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10878_ (.A1(_03112_),
    .A2(_03115_),
    .Z(_03129_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10879_ (.A1(_03128_),
    .A2(_02890_),
    .B(_03129_),
    .ZN(_03130_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10880_ (.I(_03088_),
    .Z(_03131_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10881_ (.A1(_03131_),
    .A2(_02940_),
    .ZN(_03132_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10882_ (.I0(_03130_),
    .I1(_03129_),
    .S(_03132_),
    .Z(_03133_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10883_ (.A1(_03127_),
    .A2(_03133_),
    .Z(_03134_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _10884_ (.A1(_03126_),
    .A2(_03134_),
    .Z(_03135_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _10885_ (.A1(_03125_),
    .A2(_03135_),
    .ZN(_03136_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10886_ (.A1(\channels.sample3[10] ),
    .A2(_03105_),
    .ZN(_03137_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10887_ (.A1(_03054_),
    .A2(_03136_),
    .B(_03137_),
    .ZN(_00281_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10888_ (.I(_02358_),
    .Z(_03138_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10889_ (.A1(_03127_),
    .A2(_03130_),
    .B(_03132_),
    .ZN(_03139_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10890_ (.A1(_03126_),
    .A2(_03134_),
    .ZN(_03140_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _10891_ (.A1(_03125_),
    .A2(_03135_),
    .B(_03139_),
    .C(_03140_),
    .ZN(_03141_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10892_ (.A1(_02056_),
    .A2(_03105_),
    .ZN(_03142_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10893_ (.A1(_03138_),
    .A2(_03141_),
    .B(_03142_),
    .ZN(_00282_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10894_ (.I(_01104_),
    .Z(_03143_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10895_ (.A1(\channels.sample2[0] ),
    .A2(_03143_),
    .ZN(_03144_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10896_ (.A1(_02366_),
    .A2(_02783_),
    .B(_03144_),
    .ZN(_00283_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10897_ (.A1(\channels.sample2[1] ),
    .A2(_03143_),
    .ZN(_03145_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10898_ (.A1(_02366_),
    .A2(_02831_),
    .B(_03145_),
    .ZN(_00284_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10899_ (.A1(\channels.sample2[2] ),
    .A2(_03143_),
    .ZN(_03146_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10900_ (.A1(_02366_),
    .A2(_02880_),
    .B(_03146_),
    .ZN(_00285_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10901_ (.I(_02365_),
    .Z(_03147_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10902_ (.A1(\channels.sample2[3] ),
    .A2(_03143_),
    .ZN(_03148_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10903_ (.A1(_03147_),
    .A2(_02932_),
    .B(_03148_),
    .ZN(_00286_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10904_ (.I(_01103_),
    .Z(_03149_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10905_ (.I(_03149_),
    .Z(_03150_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10906_ (.A1(\channels.sample2[4] ),
    .A2(_03150_),
    .ZN(_03151_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10907_ (.A1(_03147_),
    .A2(_02973_),
    .B(_03151_),
    .ZN(_00287_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10908_ (.A1(\channels.sample2[5] ),
    .A2(_03150_),
    .ZN(_03152_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10909_ (.A1(_03147_),
    .A2(_03013_),
    .B(_03152_),
    .ZN(_00288_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10910_ (.A1(\channels.sample2[6] ),
    .A2(_03150_),
    .ZN(_03153_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10911_ (.A1(_03147_),
    .A2(_03052_),
    .B(_03153_),
    .ZN(_00289_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10912_ (.I(_02365_),
    .Z(_03154_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10913_ (.A1(\channels.sample2[7] ),
    .A2(_03150_),
    .ZN(_03155_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10914_ (.A1(_03154_),
    .A2(_03080_),
    .B(_03155_),
    .ZN(_00290_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10915_ (.I(_03149_),
    .Z(_03156_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10916_ (.A1(\channels.sample2[8] ),
    .A2(_03156_),
    .ZN(_03157_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10917_ (.A1(_03154_),
    .A2(_03104_),
    .B(_03157_),
    .ZN(_00291_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10918_ (.A1(\channels.sample2[9] ),
    .A2(_03156_),
    .ZN(_03158_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10919_ (.A1(_03154_),
    .A2(_03122_),
    .B(_03158_),
    .ZN(_00292_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10920_ (.A1(\channels.sample2[10] ),
    .A2(_03156_),
    .ZN(_03159_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10921_ (.A1(_03154_),
    .A2(_03136_),
    .B(_03159_),
    .ZN(_00293_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10922_ (.I(_02365_),
    .Z(_03160_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10923_ (.A1(\channels.sample2[11] ),
    .A2(_03156_),
    .ZN(_03161_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10924_ (.A1(_03160_),
    .A2(_03141_),
    .B(_03161_),
    .ZN(_00294_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10925_ (.I(_01321_),
    .Z(_03162_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10926_ (.A1(\channels.sample1[0] ),
    .A2(_01560_),
    .ZN(_03163_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10927_ (.A1(_03162_),
    .A2(_02783_),
    .B(_03163_),
    .ZN(_00295_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10928_ (.I(_01460_),
    .Z(_03164_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10929_ (.A1(\channels.sample1[1] ),
    .A2(_03164_),
    .ZN(_03165_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10930_ (.A1(_03162_),
    .A2(_02831_),
    .B(_03165_),
    .ZN(_00296_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10931_ (.A1(\channels.sample1[2] ),
    .A2(_03164_),
    .ZN(_03166_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10932_ (.A1(_03162_),
    .A2(_02880_),
    .B(_03166_),
    .ZN(_00297_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10933_ (.A1(\channels.sample1[3] ),
    .A2(_03164_),
    .ZN(_03167_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10934_ (.A1(_03162_),
    .A2(_02932_),
    .B(_03167_),
    .ZN(_00298_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10935_ (.I(_01320_),
    .Z(_03168_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10936_ (.A1(\channels.sample1[4] ),
    .A2(_03164_),
    .ZN(_03169_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10937_ (.A1(_03168_),
    .A2(_02973_),
    .B(_03169_),
    .ZN(_00299_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10938_ (.I(_01460_),
    .Z(_03170_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10939_ (.A1(\channels.sample1[5] ),
    .A2(_03170_),
    .ZN(_03171_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10940_ (.A1(_03168_),
    .A2(_03013_),
    .B(_03171_),
    .ZN(_00300_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10941_ (.A1(\channels.sample1[6] ),
    .A2(_03170_),
    .ZN(_03172_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10942_ (.A1(_03168_),
    .A2(_03052_),
    .B(_03172_),
    .ZN(_00301_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10943_ (.A1(\channels.sample1[7] ),
    .A2(_03170_),
    .ZN(_03173_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10944_ (.A1(_03168_),
    .A2(_03080_),
    .B(_03173_),
    .ZN(_00302_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10945_ (.I(_01320_),
    .Z(_03174_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10946_ (.A1(\channels.sample1[8] ),
    .A2(_03170_),
    .ZN(_03175_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10947_ (.A1(_03174_),
    .A2(_03104_),
    .B(_03175_),
    .ZN(_00303_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10948_ (.A1(\channels.sample1[9] ),
    .A2(_01261_),
    .ZN(_03176_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10949_ (.A1(_03174_),
    .A2(_03122_),
    .B(_03176_),
    .ZN(_00304_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10950_ (.A1(\channels.sample1[10] ),
    .A2(_01261_),
    .ZN(_03177_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10951_ (.A1(_03174_),
    .A2(_03136_),
    .B(_03177_),
    .ZN(_00305_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10952_ (.A1(\channels.sample1[11] ),
    .A2(_01261_),
    .ZN(_03178_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10953_ (.A1(_03174_),
    .A2(_03141_),
    .B(_03178_),
    .ZN(_00306_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10954_ (.I(\filters.sample_filtered[0] ),
    .ZN(_03179_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _10955_ (.I(\filters.filter_step[2] ),
    .ZN(_03180_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _10956_ (.I(\filters.filter_step[1] ),
    .Z(_03181_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _10957_ (.I(_03181_),
    .Z(_03182_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _10958_ (.I(\filters.filter_step[0] ),
    .ZN(_03183_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _10959_ (.A1(_03180_),
    .A2(_03182_),
    .A3(_03183_),
    .ZN(_03184_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10960_ (.I(_03184_),
    .Z(_03185_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10961_ (.I(_03185_),
    .Z(_03186_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10962_ (.I(_03186_),
    .Z(_03187_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10963_ (.I(_03187_),
    .Z(_03188_));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _10964_ (.I(\filters.filter_step[2] ),
    .Z(_03189_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _10965_ (.I(_03189_),
    .Z(_03190_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _10966_ (.I(_03190_),
    .Z(_03191_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _10967_ (.I(\filters.filter_step[1] ),
    .ZN(_03192_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _10968_ (.I(_03192_),
    .Z(_03193_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _10969_ (.I(_03193_),
    .Z(_03194_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _10970_ (.I(\filters.filter_step[0] ),
    .Z(_03195_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _10971_ (.I(_03195_),
    .Z(_03196_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10972_ (.I(_03196_),
    .Z(_03197_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _10973_ (.I(\filters.band[0] ),
    .ZN(_03198_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_4 _10974_ (.A1(_03191_),
    .A2(_03194_),
    .A3(_03197_),
    .B(_03198_),
    .ZN(_03199_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10975_ (.I(_03199_),
    .Z(_03200_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10976_ (.I(_03197_),
    .Z(_03201_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10977_ (.I(_03191_),
    .Z(_03202_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _10978_ (.I(_03182_),
    .Z(_03203_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10979_ (.I(_03203_),
    .Z(_03204_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _10980_ (.A1(_03202_),
    .A2(_03204_),
    .ZN(_03205_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _10981_ (.A1(_03201_),
    .A2(_03205_),
    .ZN(_03206_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10982_ (.I(_03206_),
    .Z(_03207_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _10983_ (.A1(\filters.low[0] ),
    .A2(_03188_),
    .B(_03200_),
    .C(_03207_),
    .ZN(_03208_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10984_ (.A1(_03201_),
    .A2(_03205_),
    .Z(_03209_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10985_ (.I(_03209_),
    .Z(_03210_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10986_ (.A1(\filters.high[0] ),
    .A2(_03210_),
    .ZN(_03211_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _10987_ (.A1(_03179_),
    .A2(_03208_),
    .A3(_03211_),
    .Z(_03212_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10988_ (.A1(_03208_),
    .A2(_03211_),
    .B(_03179_),
    .ZN(_03213_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10989_ (.I(_03204_),
    .Z(_03214_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10990_ (.I(_03201_),
    .Z(_03215_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10991_ (.I(_03215_),
    .Z(_03216_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10992_ (.I(_03188_),
    .Z(_03217_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10993_ (.I(_03217_),
    .Z(_03218_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10994_ (.I(_03218_),
    .Z(_03219_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10995_ (.I(_03219_),
    .Z(_03220_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10996_ (.I(_03220_),
    .Z(_03221_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10997_ (.I(_03221_),
    .Z(_03222_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10998_ (.I(_03222_),
    .Z(_03223_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10999_ (.I(_03223_),
    .Z(_03224_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11000_ (.I(_03224_),
    .Z(_03225_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11001_ (.I(_03225_),
    .Z(_03226_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11002_ (.A1(\filters.lp ),
    .A2(_03226_),
    .ZN(_03227_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11003_ (.I(_03207_),
    .Z(_03228_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11004_ (.I(_03228_),
    .Z(_03229_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11005_ (.I(_03229_),
    .Z(_03230_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11006_ (.I(_03230_),
    .Z(_03231_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11007_ (.I(_03231_),
    .Z(_03232_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11008_ (.I(_03232_),
    .Z(_03233_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11009_ (.I(_03233_),
    .Z(_03234_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11010_ (.I(_03234_),
    .Z(_03235_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11011_ (.I(_03235_),
    .Z(_03236_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _11012_ (.A1(_03204_),
    .A2(_03215_),
    .ZN(_03237_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _11013_ (.I(_03180_),
    .Z(_03238_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _11014_ (.I(_03238_),
    .Z(_03239_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _11015_ (.A1(\filters.hp ),
    .A2(_03236_),
    .B1(_03237_),
    .B2(\filters.bp ),
    .C(_03239_),
    .ZN(_03240_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _11016_ (.A1(_01069_),
    .A2(_03227_),
    .A3(_03240_),
    .ZN(_03241_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _11017_ (.A1(_03214_),
    .A2(_03216_),
    .B(_03241_),
    .ZN(_03242_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11018_ (.I(_03242_),
    .Z(_03243_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11019_ (.I(_03241_),
    .Z(_03244_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11020_ (.I(_03244_),
    .Z(_03245_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _11021_ (.A1(_03212_),
    .A2(_03213_),
    .A3(_03243_),
    .B1(_03245_),
    .B2(_03179_),
    .ZN(_00307_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _11022_ (.I(\filters.filter_step[2] ),
    .Z(_03246_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _11023_ (.I(_03246_),
    .Z(_03247_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _11024_ (.I(_03193_),
    .Z(_03248_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _11025_ (.I(\filters.filter_step[0] ),
    .Z(_03249_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11026_ (.I(_03249_),
    .Z(_03250_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _11027_ (.I(\filters.band[1] ),
    .ZN(_03251_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _11028_ (.A1(_03247_),
    .A2(_03248_),
    .A3(_03250_),
    .B(_03251_),
    .ZN(_03252_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11029_ (.I(_03252_),
    .Z(_03253_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11030_ (.I(_03253_),
    .Z(_03254_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11031_ (.I(_03254_),
    .Z(_03255_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _11032_ (.I(_03255_),
    .Z(_03256_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _11033_ (.A1(\filters.low[1] ),
    .A2(_03187_),
    .B(_03256_),
    .C(_03206_),
    .ZN(_03257_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11034_ (.A1(\filters.high[1] ),
    .A2(_03209_),
    .ZN(_03258_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11035_ (.A1(_03257_),
    .A2(_03258_),
    .ZN(_03259_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11036_ (.A1(\filters.sample_filtered[1] ),
    .A2(_03259_),
    .Z(_03260_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11037_ (.A1(_03213_),
    .A2(_03260_),
    .Z(_03261_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11038_ (.A1(_03213_),
    .A2(_03260_),
    .ZN(_03262_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _11039_ (.I(\filters.sample_filtered[1] ),
    .ZN(_03263_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _11040_ (.A1(_03243_),
    .A2(_03261_),
    .A3(_03262_),
    .B1(_03245_),
    .B2(_03263_),
    .ZN(_00308_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11041_ (.I(\filters.sample_filtered[2] ),
    .ZN(_03264_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11042_ (.I(_03244_),
    .Z(_03265_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11043_ (.I(_03242_),
    .Z(_03266_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11044_ (.A1(_03257_),
    .A2(_03258_),
    .B(_03263_),
    .ZN(_03267_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11045_ (.I(\filters.low[2] ),
    .Z(_03268_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _11046_ (.I(\filters.band[2] ),
    .ZN(_03269_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_4 _11047_ (.A1(_03190_),
    .A2(_03193_),
    .A3(_03196_),
    .B(_03269_),
    .ZN(_03270_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11048_ (.I(_03270_),
    .Z(_03271_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11049_ (.I(_03271_),
    .Z(_03272_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11050_ (.I(_03272_),
    .Z(_03273_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _11051_ (.A1(_03268_),
    .A2(_03188_),
    .B(_03273_),
    .C(_03206_),
    .ZN(_03274_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11052_ (.A1(\filters.high[2] ),
    .A2(_03209_),
    .ZN(_03275_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11053_ (.A1(_03274_),
    .A2(_03275_),
    .ZN(_03276_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11054_ (.A1(\filters.sample_filtered[2] ),
    .A2(_03276_),
    .Z(_03277_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11055_ (.A1(_03267_),
    .A2(_03261_),
    .B(_03277_),
    .ZN(_03278_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _11056_ (.A1(_03267_),
    .A2(_03261_),
    .A3(_03277_),
    .Z(_03279_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11057_ (.A1(_03278_),
    .A2(_03279_),
    .ZN(_03280_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _11058_ (.A1(_03264_),
    .A2(_03265_),
    .B1(_03266_),
    .B2(_03280_),
    .ZN(_00309_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11059_ (.I(\filters.sample_filtered[3] ),
    .ZN(_03281_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11060_ (.I(\filters.low[3] ),
    .Z(_03282_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _11061_ (.I(_03192_),
    .Z(_03283_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _11062_ (.I(\filters.band[3] ),
    .ZN(_03284_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_4 _11063_ (.A1(_03246_),
    .A2(_03283_),
    .A3(_03249_),
    .B(_03284_),
    .ZN(_03285_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11064_ (.I(_03285_),
    .Z(_03286_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11065_ (.I(net63),
    .Z(_03287_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11066_ (.I(_03287_),
    .Z(_03288_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11067_ (.A1(_03282_),
    .A2(_03188_),
    .B(_03288_),
    .C(_03206_),
    .ZN(_03289_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11068_ (.A1(\filters.high[3] ),
    .A2(_03210_),
    .ZN(_03290_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11069_ (.A1(_03289_),
    .A2(_03290_),
    .ZN(_03291_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11070_ (.A1(\filters.sample_filtered[3] ),
    .A2(_03291_),
    .Z(_03292_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11071_ (.I(_03292_),
    .ZN(_03293_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11072_ (.A1(\filters.sample_filtered[2] ),
    .A2(_03276_),
    .ZN(_03294_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11073_ (.A1(_03294_),
    .A2(_03278_),
    .ZN(_03295_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11074_ (.A1(_03293_),
    .A2(_03295_),
    .Z(_03296_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _11075_ (.A1(_03281_),
    .A2(_03265_),
    .B1(_03266_),
    .B2(_03296_),
    .ZN(_00310_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11076_ (.I(\filters.sample_filtered[4] ),
    .ZN(_03297_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _11077_ (.I(\filters.high[4] ),
    .ZN(_03298_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_3 _11078_ (.I(\filters.band[4] ),
    .ZN(_03299_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_4 _11079_ (.A1(_03246_),
    .A2(_03283_),
    .A3(_03249_),
    .B(_03299_),
    .ZN(_03300_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11080_ (.I(_03300_),
    .Z(_03301_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11081_ (.I(_03301_),
    .Z(_03302_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11082_ (.A1(\filters.low[4] ),
    .A2(_03217_),
    .B(_03302_),
    .C(_03207_),
    .ZN(_03303_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _11083_ (.A1(_03298_),
    .A2(_03207_),
    .B(_03303_),
    .ZN(_03304_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11084_ (.A1(\filters.sample_filtered[4] ),
    .A2(_03304_),
    .Z(_03305_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11085_ (.A1(_03294_),
    .A2(_03278_),
    .B(_03293_),
    .ZN(_03306_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _11086_ (.A1(\filters.sample_filtered[3] ),
    .A2(_03291_),
    .B(_03306_),
    .ZN(_03307_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11087_ (.A1(_03305_),
    .A2(_03307_),
    .Z(_03308_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _11088_ (.A1(_03297_),
    .A2(_03265_),
    .B1(_03266_),
    .B2(_03308_),
    .ZN(_00311_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _11089_ (.I(\filters.sample_filtered[5] ),
    .ZN(_03309_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11090_ (.I(\filters.low[5] ),
    .Z(_03310_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _11091_ (.I(_03189_),
    .Z(_03311_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _11092_ (.I(_03283_),
    .Z(_03312_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _11093_ (.I(_03195_),
    .Z(_03313_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _11094_ (.I(\filters.band[5] ),
    .ZN(_03314_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_4 _11095_ (.A1(_03311_),
    .A2(_03312_),
    .A3(_03313_),
    .B(_03314_),
    .ZN(_03315_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11096_ (.I(_03315_),
    .Z(_03316_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11097_ (.I(_03316_),
    .Z(_03317_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _11098_ (.A1(_03310_),
    .A2(_03217_),
    .B(_03317_),
    .C(_03228_),
    .ZN(_03318_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11099_ (.A1(\filters.high[5] ),
    .A2(_03210_),
    .ZN(_03319_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11100_ (.A1(_03318_),
    .A2(_03319_),
    .ZN(_03320_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11101_ (.A1(\filters.sample_filtered[5] ),
    .A2(_03320_),
    .Z(_03321_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11102_ (.I(_03305_),
    .ZN(_03322_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11103_ (.A1(\filters.sample_filtered[4] ),
    .A2(_03304_),
    .ZN(_03323_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _11104_ (.A1(_03322_),
    .A2(_03307_),
    .B(_03323_),
    .ZN(_03324_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _11105_ (.A1(_03321_),
    .A2(_03324_),
    .ZN(_03325_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _11106_ (.A1(_03309_),
    .A2(_03265_),
    .B1(_03266_),
    .B2(_03325_),
    .ZN(_00312_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11107_ (.I(\filters.sample_filtered[6] ),
    .ZN(_03326_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11108_ (.I(_03244_),
    .Z(_03327_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11109_ (.I(_03242_),
    .Z(_03328_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11110_ (.I(\filters.low[6] ),
    .Z(_03329_));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 _11111_ (.I(\filters.band[6] ),
    .ZN(_03330_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _11112_ (.A1(_03247_),
    .A2(_03248_),
    .A3(_03250_),
    .B(_03330_),
    .ZN(_03331_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11113_ (.I(_03331_),
    .Z(_03332_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11114_ (.I(_03332_),
    .Z(_03333_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _11115_ (.A1(_03329_),
    .A2(_03218_),
    .B(_03333_),
    .C(_03228_),
    .ZN(_03334_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11116_ (.I(_03210_),
    .Z(_03335_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11117_ (.A1(\filters.high[6] ),
    .A2(_03335_),
    .ZN(_03336_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _11118_ (.A1(_03334_),
    .A2(_03336_),
    .ZN(_03337_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11119_ (.A1(\filters.sample_filtered[6] ),
    .A2(_03337_),
    .Z(_03338_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11120_ (.A1(_03318_),
    .A2(_03319_),
    .B(_03309_),
    .ZN(_03339_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _11121_ (.A1(_03321_),
    .A2(_03324_),
    .B(_03339_),
    .ZN(_03340_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11122_ (.A1(_03338_),
    .A2(_03340_),
    .Z(_03341_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _11123_ (.A1(_03326_),
    .A2(_03327_),
    .B1(_03328_),
    .B2(_03341_),
    .ZN(_00313_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11124_ (.I(\filters.sample_filtered[7] ),
    .ZN(_03342_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _11125_ (.I(\filters.high[7] ),
    .ZN(_03343_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11126_ (.I(_03228_),
    .Z(_03344_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11127_ (.I(\filters.low[7] ),
    .Z(_03345_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11128_ (.I(_03218_),
    .Z(_03346_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _11129_ (.I(\filters.band[7] ),
    .ZN(_03347_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_4 _11130_ (.A1(_03191_),
    .A2(_03248_),
    .A3(_03197_),
    .B(_03347_),
    .ZN(_03348_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11131_ (.I(_03348_),
    .Z(_03349_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _11132_ (.I(_03349_),
    .Z(_03350_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _11133_ (.A1(_03345_),
    .A2(_03346_),
    .B(_03350_),
    .C(_03229_),
    .ZN(_03351_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _11134_ (.A1(_03343_),
    .A2(_03344_),
    .B(_03351_),
    .ZN(_03352_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11135_ (.A1(\filters.sample_filtered[7] ),
    .A2(_03352_),
    .Z(_03353_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11136_ (.I(_03338_),
    .ZN(_03354_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11137_ (.A1(_03354_),
    .A2(_03340_),
    .ZN(_03355_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _11138_ (.A1(\filters.sample_filtered[6] ),
    .A2(_03337_),
    .B(_03355_),
    .ZN(_03356_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11139_ (.A1(_03353_),
    .A2(_03356_),
    .Z(_03357_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _11140_ (.A1(_03342_),
    .A2(_03327_),
    .B1(_03328_),
    .B2(_03357_),
    .ZN(_00314_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11141_ (.I(\filters.sample_filtered[8] ),
    .ZN(_03358_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _11142_ (.I(\filters.high[8] ),
    .ZN(_03359_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11143_ (.I(\filters.low[8] ),
    .Z(_03360_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _11144_ (.I(\filters.band[8] ),
    .ZN(_03361_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_4 _11145_ (.A1(_03191_),
    .A2(_03248_),
    .A3(_03197_),
    .B(_03361_),
    .ZN(_03362_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _11146_ (.I(_03362_),
    .Z(_03363_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _11147_ (.I(_03363_),
    .Z(_03364_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _11148_ (.A1(_03360_),
    .A2(_03220_),
    .B(_03364_),
    .C(_03344_),
    .ZN(_03365_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _11149_ (.A1(_03359_),
    .A2(_03230_),
    .B(_03365_),
    .ZN(_03366_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11150_ (.A1(\filters.sample_filtered[8] ),
    .A2(_03366_),
    .Z(_03367_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11151_ (.I(_03353_),
    .ZN(_03368_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11152_ (.A1(_03368_),
    .A2(_03356_),
    .ZN(_03369_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11153_ (.A1(\filters.sample_filtered[7] ),
    .A2(_03352_),
    .B(_03369_),
    .ZN(_03370_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11154_ (.A1(_03367_),
    .A2(_03370_),
    .Z(_03371_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _11155_ (.A1(_03358_),
    .A2(_03327_),
    .B1(_03328_),
    .B2(_03371_),
    .ZN(_00315_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11156_ (.I(\filters.sample_filtered[9] ),
    .ZN(_03372_));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 _11157_ (.I(\filters.high[9] ),
    .ZN(_03373_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11158_ (.I(\filters.low[9] ),
    .Z(_03374_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11159_ (.I(_03217_),
    .Z(_03375_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11160_ (.I(_03375_),
    .Z(_03376_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11161_ (.I(_03376_),
    .Z(_03377_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11162_ (.I(_03377_),
    .Z(_03378_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _11163_ (.I(_03283_),
    .Z(_03379_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _11164_ (.I(\filters.band[9] ),
    .ZN(_03380_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_4 _11165_ (.A1(_03247_),
    .A2(_03379_),
    .A3(_03250_),
    .B(_03380_),
    .ZN(_03381_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11166_ (.I(_03381_),
    .Z(_03382_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11167_ (.I(_03382_),
    .Z(_03383_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _11168_ (.A1(_03374_),
    .A2(_03378_),
    .B(_03383_),
    .C(_03230_),
    .ZN(_03384_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _11169_ (.A1(_03373_),
    .A2(_03231_),
    .B(_03384_),
    .ZN(_03385_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11170_ (.A1(\filters.sample_filtered[9] ),
    .A2(_03385_),
    .Z(_03386_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11171_ (.I(_03367_),
    .ZN(_03387_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11172_ (.A1(_03387_),
    .A2(_03370_),
    .ZN(_03388_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11173_ (.A1(\filters.sample_filtered[8] ),
    .A2(_03366_),
    .B(_03388_),
    .ZN(_03389_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11174_ (.A1(_03386_),
    .A2(_03389_),
    .Z(_03390_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _11175_ (.A1(_03372_),
    .A2(_03327_),
    .B1(_03328_),
    .B2(_03390_),
    .ZN(_00316_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _11176_ (.I(\filters.sample_filtered[10] ),
    .ZN(_03391_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11177_ (.I(_03244_),
    .Z(_03392_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11178_ (.I(_03242_),
    .Z(_03393_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11179_ (.I(\filters.low[10] ),
    .Z(_03394_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11180_ (.I(_03221_),
    .Z(_03395_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _11181_ (.I(\filters.band[10] ),
    .ZN(_03396_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_4 _11182_ (.A1(_03247_),
    .A2(_03379_),
    .A3(_03250_),
    .B(_03396_),
    .ZN(_03397_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11183_ (.I(_03397_),
    .Z(_03398_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11184_ (.A1(_03394_),
    .A2(_03395_),
    .B(_03398_),
    .C(_03232_),
    .ZN(_03399_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11185_ (.I(_03335_),
    .Z(_03400_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11186_ (.I(_03400_),
    .Z(_03401_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11187_ (.A1(\filters.high[10] ),
    .A2(_03401_),
    .ZN(_03402_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11188_ (.A1(_03399_),
    .A2(_03402_),
    .ZN(_03403_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11189_ (.A1(\filters.sample_filtered[10] ),
    .A2(_03403_),
    .Z(_03404_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11190_ (.I(_03386_),
    .ZN(_03405_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11191_ (.A1(_03405_),
    .A2(_03389_),
    .ZN(_03406_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11192_ (.A1(\filters.sample_filtered[9] ),
    .A2(_03385_),
    .B(_03406_),
    .ZN(_03407_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11193_ (.A1(_03404_),
    .A2(_03407_),
    .Z(_03408_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _11194_ (.A1(_03391_),
    .A2(_03392_),
    .B1(_03393_),
    .B2(_03408_),
    .ZN(_00317_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11195_ (.I(\filters.sample_filtered[11] ),
    .ZN(_03409_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _11196_ (.I(\filters.high[11] ),
    .ZN(_03410_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11197_ (.I(\filters.low[11] ),
    .Z(_03411_));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 _11198_ (.I(\filters.band[11] ),
    .ZN(_03412_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_4 _11199_ (.A1(_03311_),
    .A2(_03379_),
    .A3(_03313_),
    .B(_03412_),
    .ZN(_03413_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _11200_ (.A1(_03411_),
    .A2(_03223_),
    .B(_03413_),
    .C(_03233_),
    .ZN(_03414_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _11201_ (.A1(_03410_),
    .A2(_03233_),
    .B(_03414_),
    .ZN(_03415_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11202_ (.A1(\filters.sample_filtered[11] ),
    .A2(_03415_),
    .Z(_03416_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11203_ (.I(_03404_),
    .ZN(_03417_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11204_ (.A1(_03417_),
    .A2(_03407_),
    .ZN(_03418_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11205_ (.A1(\filters.sample_filtered[10] ),
    .A2(_03403_),
    .B(_03418_),
    .ZN(_03419_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11206_ (.A1(_03416_),
    .A2(_03419_),
    .Z(_03420_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _11207_ (.A1(_03409_),
    .A2(_03392_),
    .B1(_03393_),
    .B2(_03420_),
    .ZN(_00318_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11208_ (.I(\filters.sample_filtered[12] ),
    .ZN(_03421_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11209_ (.I(\filters.low[12] ),
    .Z(_03422_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _11210_ (.I(\filters.band[12] ),
    .ZN(_03423_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11211_ (.I(_03395_),
    .Z(_03424_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11212_ (.A1(_03423_),
    .A2(_03424_),
    .ZN(_03425_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _11213_ (.A1(_03422_),
    .A2(_03224_),
    .B(_03425_),
    .C(_03234_),
    .ZN(_03426_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11214_ (.I(_03401_),
    .Z(_03427_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11215_ (.I(_03427_),
    .Z(_03428_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11216_ (.A1(\filters.high[12] ),
    .A2(_03428_),
    .ZN(_03429_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11217_ (.A1(_03426_),
    .A2(_03429_),
    .ZN(_03430_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11218_ (.A1(\filters.sample_filtered[12] ),
    .A2(_03430_),
    .Z(_03431_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11219_ (.I(_03416_),
    .ZN(_03432_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11220_ (.A1(_03432_),
    .A2(_03419_),
    .ZN(_03433_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11221_ (.A1(\filters.sample_filtered[11] ),
    .A2(_03415_),
    .B(_03433_),
    .ZN(_03434_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11222_ (.A1(_03431_),
    .A2(_03434_),
    .Z(_03435_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _11223_ (.A1(_03421_),
    .A2(_03392_),
    .B1(_03393_),
    .B2(_03435_),
    .ZN(_00319_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11224_ (.A1(_03426_),
    .A2(_03429_),
    .B(_03421_),
    .ZN(_03436_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11225_ (.I(_03431_),
    .ZN(_03437_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11226_ (.A1(_03437_),
    .A2(_03434_),
    .ZN(_03438_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11227_ (.I(\filters.low[13] ),
    .Z(_03439_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _11228_ (.I(\filters.band[13] ),
    .ZN(_03440_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11229_ (.A1(_03440_),
    .A2(_03224_),
    .ZN(_03441_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11230_ (.A1(_03439_),
    .A2(_03225_),
    .B(_03441_),
    .ZN(_03442_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11231_ (.A1(\filters.high[13] ),
    .A2(_03235_),
    .ZN(_03443_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _11232_ (.A1(_03235_),
    .A2(_03442_),
    .B(_03443_),
    .ZN(_03444_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11233_ (.A1(\filters.sample_filtered[13] ),
    .A2(_03444_),
    .Z(_03445_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _11234_ (.A1(_03436_),
    .A2(_03438_),
    .A3(_03445_),
    .ZN(_03446_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11235_ (.I(_03445_),
    .ZN(_03447_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11236_ (.A1(_03436_),
    .A2(_03438_),
    .ZN(_03448_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11237_ (.A1(_03447_),
    .A2(_03448_),
    .ZN(_03449_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11238_ (.I(\filters.sample_filtered[13] ),
    .Z(_03450_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11239_ (.I(_03450_),
    .ZN(_03451_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _11240_ (.A1(_03243_),
    .A2(_03446_),
    .A3(_03449_),
    .B1(_03245_),
    .B2(_03451_),
    .ZN(_00320_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11241_ (.I(\filters.sample_filtered[14] ),
    .Z(_03452_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11242_ (.I(_03452_),
    .ZN(_03453_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11243_ (.A1(_03450_),
    .A2(_03444_),
    .B(_03449_),
    .ZN(_03454_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11244_ (.I(\filters.low[14] ),
    .Z(_03455_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _11245_ (.I(\filters.band[14] ),
    .ZN(_03456_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11246_ (.A1(_03456_),
    .A2(_03225_),
    .ZN(_03457_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11247_ (.A1(_03455_),
    .A2(_03226_),
    .B(_03457_),
    .ZN(_03458_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11248_ (.A1(\filters.high[14] ),
    .A2(_03235_),
    .ZN(_03459_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _11249_ (.A1(_03236_),
    .A2(_03458_),
    .B(_03459_),
    .ZN(_03460_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11250_ (.A1(_03452_),
    .A2(_03460_),
    .Z(_03461_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11251_ (.A1(_03454_),
    .A2(_03461_),
    .Z(_03462_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _11252_ (.A1(_03453_),
    .A2(_03392_),
    .B1(_03393_),
    .B2(_03462_),
    .ZN(_00321_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11253_ (.I(_03461_),
    .ZN(_03463_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11254_ (.A1(_03454_),
    .A2(_03463_),
    .ZN(_03464_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11255_ (.A1(_03452_),
    .A2(_03460_),
    .B(_03464_),
    .ZN(_03465_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11256_ (.I(\filters.sample_filtered[15] ),
    .ZN(_03466_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11257_ (.I(\filters.high[15] ),
    .ZN(_03467_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11258_ (.I(\filters.low[15] ),
    .Z(_03468_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11259_ (.A1(_03468_),
    .A2(_03226_),
    .ZN(_03469_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _11260_ (.A1(_03202_),
    .A2(_03194_),
    .A3(_03201_),
    .ZN(_03470_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11261_ (.I(_03470_),
    .Z(_03471_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11262_ (.I(_03471_),
    .Z(_03472_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11263_ (.I(_03472_),
    .Z(_03473_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11264_ (.I(_03473_),
    .Z(_03474_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11265_ (.I(_03474_),
    .Z(_03475_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11266_ (.I(_03475_),
    .Z(_03476_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11267_ (.I(_03476_),
    .Z(_03477_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11268_ (.A1(\filters.band[15] ),
    .A2(_03477_),
    .B(_03236_),
    .ZN(_03478_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _11269_ (.A1(_03467_),
    .A2(_03236_),
    .B1(_03469_),
    .B2(_03478_),
    .ZN(_03479_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11270_ (.A1(_03466_),
    .A2(_03479_),
    .Z(_03480_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11271_ (.A1(_03465_),
    .A2(_03480_),
    .Z(_03481_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11272_ (.A1(_03465_),
    .A2(_03480_),
    .ZN(_03482_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _11273_ (.A1(_03243_),
    .A2(_03481_),
    .A3(_03482_),
    .B1(_03245_),
    .B2(_03466_),
    .ZN(_00322_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11274_ (.A1(_02088_),
    .A2(_01849_),
    .Z(_03483_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11275_ (.I(_03483_),
    .Z(_03484_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11276_ (.I(_02334_),
    .Z(_03485_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11277_ (.A1(\filters.cutoff_lut[6] ),
    .A2(_03484_),
    .B(_03485_),
    .ZN(_03486_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11278_ (.A1(_02308_),
    .A2(_03484_),
    .B(_03486_),
    .ZN(_00323_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11279_ (.A1(\filters.cutoff_lut[7] ),
    .A2(_03483_),
    .B(_03485_),
    .ZN(_03487_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11280_ (.A1(_02314_),
    .A2(_03484_),
    .B(_03487_),
    .ZN(_00324_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11281_ (.A1(\filters.cutoff_lut[8] ),
    .A2(_03483_),
    .B(_03485_),
    .ZN(_03488_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11282_ (.A1(_02316_),
    .A2(_03484_),
    .B(_03488_),
    .ZN(_00325_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11283_ (.I(\tt_um_rejunity_sn76489.control_tone_freq[0][0] ),
    .ZN(_03489_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11284_ (.I(net14),
    .Z(_03490_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11285_ (.I(net13),
    .Z(_03491_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11286_ (.I(net12),
    .Z(_03492_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11287_ (.A1(_00999_),
    .A2(_01003_),
    .ZN(_03493_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _11288_ (.A1(_01824_),
    .A2(_01093_),
    .A3(_01831_),
    .A4(_03493_),
    .ZN(_03494_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _11289_ (.A1(net15),
    .A2(_03494_),
    .ZN(_03495_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11290_ (.I(_03495_),
    .Z(_03496_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _11291_ (.A1(_03490_),
    .A2(_03491_),
    .A3(_03492_),
    .A4(_03496_),
    .ZN(_03497_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11292_ (.I(_03497_),
    .Z(_03498_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11293_ (.I(net8),
    .Z(_03499_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11294_ (.I(_03497_),
    .Z(_03500_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11295_ (.A1(_03499_),
    .A2(_03500_),
    .ZN(_03501_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11296_ (.A1(_03489_),
    .A2(_03498_),
    .B(_03501_),
    .C(_02273_),
    .ZN(_00326_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11297_ (.A1(\tt_um_rejunity_sn76489.control_tone_freq[0][1] ),
    .A2(_03500_),
    .B(_03485_),
    .ZN(_03502_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11298_ (.A1(_02314_),
    .A2(_03498_),
    .B(_03502_),
    .ZN(_00327_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11299_ (.I(_02334_),
    .Z(_03503_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11300_ (.A1(\tt_um_rejunity_sn76489.control_tone_freq[0][2] ),
    .A2(_03500_),
    .B(_03503_),
    .ZN(_03504_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11301_ (.A1(_02316_),
    .A2(_03498_),
    .B(_03504_),
    .ZN(_00328_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11302_ (.A1(\tt_um_rejunity_sn76489.control_tone_freq[0][3] ),
    .A2(_03500_),
    .B(_03503_),
    .ZN(_03505_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11303_ (.A1(_02299_),
    .A2(_03498_),
    .B(_03505_),
    .ZN(_00329_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11304_ (.I(\tt_um_rejunity_sn76489.control_tone_freq[2][0] ),
    .ZN(_03506_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _11305_ (.A1(_01812_),
    .A2(_03491_),
    .A3(_03492_),
    .A4(_03495_),
    .ZN(_03507_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11306_ (.I(_03507_),
    .Z(_03508_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11307_ (.I(_03507_),
    .Z(_03509_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11308_ (.A1(_03499_),
    .A2(_03509_),
    .ZN(_03510_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11309_ (.A1(_03506_),
    .A2(_03508_),
    .B(_03510_),
    .C(_02273_),
    .ZN(_00330_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11310_ (.I(_02184_),
    .Z(_03511_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11311_ (.A1(\tt_um_rejunity_sn76489.control_tone_freq[2][1] ),
    .A2(_03509_),
    .B(_03503_),
    .ZN(_03512_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11312_ (.A1(_03511_),
    .A2(_03508_),
    .B(_03512_),
    .ZN(_00331_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11313_ (.I(_02187_),
    .Z(_03513_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11314_ (.A1(\tt_um_rejunity_sn76489.control_tone_freq[2][2] ),
    .A2(_03509_),
    .B(_03503_),
    .ZN(_03514_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11315_ (.A1(_03513_),
    .A2(_03508_),
    .B(_03514_),
    .ZN(_00332_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11316_ (.I(_02298_),
    .Z(_03515_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11317_ (.I(_02333_),
    .Z(_03516_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11318_ (.I(_03516_),
    .Z(_03517_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11319_ (.A1(\tt_um_rejunity_sn76489.control_tone_freq[2][3] ),
    .A2(_03509_),
    .B(_03517_),
    .ZN(_03518_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11320_ (.A1(_03515_),
    .A2(_03508_),
    .B(_03518_),
    .ZN(_00333_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _11321_ (.A1(_01805_),
    .A2(_03492_),
    .ZN(_03519_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11322_ (.A1(_01811_),
    .A2(_03495_),
    .ZN(_03520_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11323_ (.A1(_03519_),
    .A2(_03520_),
    .Z(_03521_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11324_ (.I(_03521_),
    .Z(_03522_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11325_ (.I(_03521_),
    .Z(_03523_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11326_ (.A1(_01740_),
    .A2(_03523_),
    .ZN(_03524_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11327_ (.A1(\tt_um_rejunity_sn76489.control_tone_freq[1][0] ),
    .A2(_03522_),
    .B(_03524_),
    .ZN(_03525_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11328_ (.A1(_02103_),
    .A2(_03525_),
    .ZN(_00334_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11329_ (.A1(\tt_um_rejunity_sn76489.control_tone_freq[1][1] ),
    .A2(_03523_),
    .B(_03517_),
    .ZN(_03526_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11330_ (.A1(_03511_),
    .A2(_03522_),
    .B(_03526_),
    .ZN(_00335_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11331_ (.A1(\tt_um_rejunity_sn76489.control_tone_freq[1][2] ),
    .A2(_03523_),
    .B(_03517_),
    .ZN(_03527_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11332_ (.A1(_03513_),
    .A2(_03522_),
    .B(_03527_),
    .ZN(_00336_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11333_ (.A1(\tt_um_rejunity_sn76489.control_tone_freq[1][3] ),
    .A2(_03523_),
    .B(_03517_),
    .ZN(_03528_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11334_ (.A1(_03515_),
    .A2(_03522_),
    .B(_03528_),
    .ZN(_00337_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _11335_ (.I0(\channels.adsr_state[0][0] ),
    .I1(\channels.adsr_state[1][0] ),
    .I2(\channels.adsr_state[2][0] ),
    .I3(\channels.adsr_state[3][0] ),
    .S0(_01146_),
    .S1(_01160_),
    .Z(_03529_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11336_ (.I(_03529_),
    .ZN(_03530_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _11337_ (.I0(\channels.adsr_state[0][1] ),
    .I1(\channels.adsr_state[1][1] ),
    .I2(\channels.adsr_state[2][1] ),
    .I3(\channels.adsr_state[3][1] ),
    .S0(_01147_),
    .S1(_01161_),
    .Z(_03531_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _11338_ (.A1(_03530_),
    .A2(_03531_),
    .ZN(_03532_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11339_ (.I(_03532_),
    .Z(_03533_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11340_ (.I(_03533_),
    .Z(_03534_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11341_ (.I(_02805_),
    .Z(_03535_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11342_ (.I(_02710_),
    .Z(_03536_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11343_ (.A1(_02707_),
    .A2(_02711_),
    .ZN(_03537_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11344_ (.A1(_03039_),
    .A2(_03536_),
    .A3(_03537_),
    .ZN(_03538_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11345_ (.I(_03096_),
    .Z(_03539_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11346_ (.I(_03028_),
    .Z(_03540_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11347_ (.A1(_03539_),
    .A2(_03540_),
    .ZN(_03541_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _11348_ (.A1(_03538_),
    .A2(_03541_),
    .Z(_03542_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _11349_ (.A1(_03535_),
    .A2(_03542_),
    .Z(_03543_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _11350_ (.A1(_02847_),
    .A2(_03543_),
    .ZN(_03544_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _11351_ (.A1(_01585_),
    .A2(_03534_),
    .A3(_03544_),
    .ZN(_03545_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11352_ (.A1(_03534_),
    .A2(_03544_),
    .ZN(_03546_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11353_ (.A1(\channels.ctrl_reg2[0] ),
    .A2(_01282_),
    .ZN(_03547_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11354_ (.A1(\channels.ctrl_reg3[0] ),
    .A2(_01581_),
    .B1(_01295_),
    .B2(\channels.ctrl_reg1[0] ),
    .ZN(_03548_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _11355_ (.A1(_03547_),
    .A2(_03548_),
    .ZN(_03549_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _11356_ (.A1(_03529_),
    .A2(_03531_),
    .ZN(_03550_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _11357_ (.A1(_03546_),
    .A2(_03549_),
    .A3(_03550_),
    .ZN(_03551_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _11358_ (.A1(_01254_),
    .A2(_03551_),
    .B(_01931_),
    .ZN(_03552_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11359_ (.I0(_03545_),
    .I1(\channels.adsr_state[0][0] ),
    .S(_03552_),
    .Z(_03553_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11360_ (.I(_03553_),
    .Z(_00338_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _11361_ (.A1(_01585_),
    .A2(_03529_),
    .A3(_03531_),
    .A4(_03549_),
    .ZN(_03554_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11362_ (.I0(_03554_),
    .I1(\channels.adsr_state[0][1] ),
    .S(_03552_),
    .Z(_03555_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11363_ (.I(_03555_),
    .Z(_00339_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11364_ (.I(_01088_),
    .Z(_03556_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11365_ (.I(_03556_),
    .Z(_03557_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11366_ (.I(_01084_),
    .Z(_03558_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11367_ (.A1(_01311_),
    .A2(_03557_),
    .B1(_01316_),
    .B2(_03558_),
    .ZN(_00340_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11368_ (.I(_02974_),
    .Z(_03559_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11369_ (.A1(\channels.accum[2][1] ),
    .A2(_03559_),
    .ZN(_03560_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11370_ (.A1(_03138_),
    .A2(_01333_),
    .B(_03560_),
    .ZN(_00341_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11371_ (.I(\channels.accum[2][2] ),
    .ZN(_03561_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11372_ (.A1(_03561_),
    .A2(_03557_),
    .B1(_01348_),
    .B2(_03558_),
    .ZN(_00342_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11373_ (.A1(\channels.accum[2][3] ),
    .A2(_03559_),
    .ZN(_03562_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11374_ (.A1(_03138_),
    .A2(_01359_),
    .B(_03562_),
    .ZN(_00343_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11375_ (.I(\channels.accum[2][4] ),
    .ZN(_03563_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11376_ (.A1(_03563_),
    .A2(_03557_),
    .B1(_01372_),
    .B2(_03558_),
    .ZN(_00344_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11377_ (.A1(\channels.accum[2][5] ),
    .A2(_03559_),
    .ZN(_03564_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11378_ (.A1(_03138_),
    .A2(_01381_),
    .B(_03564_),
    .ZN(_00345_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11379_ (.I(\channels.accum[2][6] ),
    .ZN(_03565_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11380_ (.A1(_03565_),
    .A2(_03557_),
    .B1(_01395_),
    .B2(_03558_),
    .ZN(_00346_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11381_ (.I(_02357_),
    .Z(_03566_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11382_ (.A1(\channels.accum[2][7] ),
    .A2(_03559_),
    .ZN(_03567_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11383_ (.A1(_03566_),
    .A2(_01406_),
    .B(_03567_),
    .ZN(_00347_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11384_ (.I(\channels.accum[2][8] ),
    .ZN(_03568_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11385_ (.I(_01089_),
    .Z(_03569_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11386_ (.I(_01240_),
    .Z(_03570_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11387_ (.A1(_03568_),
    .A2(_03569_),
    .B1(_01420_),
    .B2(_03570_),
    .ZN(_00348_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11388_ (.I(_02974_),
    .Z(_03571_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11389_ (.A1(\channels.accum[2][9] ),
    .A2(_03571_),
    .ZN(_03572_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11390_ (.A1(_03566_),
    .A2(_01433_),
    .B(_03572_),
    .ZN(_00349_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11391_ (.I(\channels.accum[2][10] ),
    .ZN(_03573_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11392_ (.A1(_03573_),
    .A2(_03569_),
    .B1(_01448_),
    .B2(_03570_),
    .ZN(_00350_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11393_ (.A1(\channels.accum[2][11] ),
    .A2(_03571_),
    .ZN(_03574_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11394_ (.A1(_03566_),
    .A2(_01459_),
    .B(_03574_),
    .ZN(_00351_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11395_ (.I(\channels.accum[2][12] ),
    .ZN(_03575_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11396_ (.A1(_03575_),
    .A2(_03569_),
    .B1(_01475_),
    .B2(_03570_),
    .ZN(_00352_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11397_ (.A1(\channels.accum[2][13] ),
    .A2(_03571_),
    .ZN(_03576_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11398_ (.A1(_03566_),
    .A2(_01487_),
    .B(_03576_),
    .ZN(_00353_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11399_ (.I(\channels.accum[2][14] ),
    .ZN(_03577_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11400_ (.A1(_03577_),
    .A2(_03569_),
    .B1(_01503_),
    .B2(_03570_),
    .ZN(_00354_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11401_ (.I(_02357_),
    .Z(_03578_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11402_ (.A1(\channels.accum[2][15] ),
    .A2(_03571_),
    .ZN(_03579_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11403_ (.A1(_03578_),
    .A2(_01515_),
    .B(_03579_),
    .ZN(_00355_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11404_ (.I(\channels.accum[2][16] ),
    .ZN(_03580_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11405_ (.I(_01089_),
    .Z(_03581_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11406_ (.I(_01240_),
    .Z(_03582_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11407_ (.A1(_03580_),
    .A2(_03581_),
    .B1(_01524_),
    .B2(_03582_),
    .ZN(_00356_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11408_ (.A1(\channels.accum[2][17] ),
    .A2(_01245_),
    .B1(_01530_),
    .B2(_01084_),
    .ZN(_03583_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11409_ (.I(_03583_),
    .ZN(_00357_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11410_ (.I(\channels.accum[2][18] ),
    .ZN(_03584_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11411_ (.A1(_03584_),
    .A2(_03581_),
    .B1(_01539_),
    .B2(_03582_),
    .ZN(_00358_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11412_ (.A1(\channels.accum[2][19] ),
    .A2(_03556_),
    .ZN(_03585_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11413_ (.A1(_03578_),
    .A2(_01545_),
    .B(_03585_),
    .ZN(_00359_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11414_ (.I(\channels.accum[2][20] ),
    .ZN(_03586_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11415_ (.A1(_03586_),
    .A2(_03581_),
    .B1(_01552_),
    .B2(_03582_),
    .ZN(_00360_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11416_ (.A1(\channels.accum[2][21] ),
    .A2(_03556_),
    .ZN(_03587_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11417_ (.A1(_03578_),
    .A2(_01559_),
    .B(_03587_),
    .ZN(_00361_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11418_ (.A1(_01564_),
    .A2(_03581_),
    .B1(_01568_),
    .B2(_03582_),
    .ZN(_00362_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11419_ (.A1(\channels.accum[2][23] ),
    .A2(_03556_),
    .ZN(_03588_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11420_ (.A1(_03578_),
    .A2(_01571_),
    .B(_03588_),
    .ZN(_00363_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11421_ (.I(\channels.accum[1][0] ),
    .ZN(_03589_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11422_ (.I(_01103_),
    .Z(_03590_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11423_ (.I(_03590_),
    .Z(_03591_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11424_ (.I(_01101_),
    .Z(_03592_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11425_ (.A1(_03589_),
    .A2(_03591_),
    .B1(_01316_),
    .B2(_03592_),
    .ZN(_00364_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11426_ (.I(_03149_),
    .Z(_03593_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11427_ (.A1(\channels.accum[1][1] ),
    .A2(_03593_),
    .ZN(_03594_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11428_ (.A1(_03160_),
    .A2(_01333_),
    .B(_03594_),
    .ZN(_00365_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11429_ (.I(\channels.accum[1][2] ),
    .ZN(_03595_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11430_ (.A1(_03595_),
    .A2(_03591_),
    .B1(_01348_),
    .B2(_03592_),
    .ZN(_00366_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11431_ (.A1(\channels.accum[1][3] ),
    .A2(_03593_),
    .ZN(_03596_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11432_ (.A1(_03160_),
    .A2(_01359_),
    .B(_03596_),
    .ZN(_00367_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11433_ (.I(\channels.accum[1][4] ),
    .ZN(_03597_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11434_ (.A1(_03597_),
    .A2(_03591_),
    .B1(_01372_),
    .B2(_03592_),
    .ZN(_00368_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11435_ (.A1(\channels.accum[1][5] ),
    .A2(_03593_),
    .ZN(_03598_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11436_ (.A1(_03160_),
    .A2(_01381_),
    .B(_03598_),
    .ZN(_00369_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11437_ (.I(\channels.accum[1][6] ),
    .ZN(_03599_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11438_ (.A1(_03599_),
    .A2(_03591_),
    .B1(_01395_),
    .B2(_03592_),
    .ZN(_00370_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11439_ (.I(_02364_),
    .Z(_03600_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11440_ (.A1(\channels.accum[1][7] ),
    .A2(_03593_),
    .ZN(_03601_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11441_ (.A1(_03600_),
    .A2(_01406_),
    .B(_03601_),
    .ZN(_00371_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11442_ (.I(\channels.accum[1][8] ),
    .ZN(_03602_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11443_ (.I(_01104_),
    .Z(_03603_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11444_ (.I(_01219_),
    .Z(_03604_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11445_ (.A1(_03602_),
    .A2(_03603_),
    .B1(_01420_),
    .B2(_03604_),
    .ZN(_00372_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11446_ (.I(_03149_),
    .Z(_03605_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11447_ (.A1(\channels.accum[1][9] ),
    .A2(_03605_),
    .ZN(_03606_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11448_ (.A1(_03600_),
    .A2(_01433_),
    .B(_03606_),
    .ZN(_00373_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11449_ (.I(\channels.accum[1][10] ),
    .ZN(_03607_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11450_ (.A1(_03607_),
    .A2(_03603_),
    .B1(_01448_),
    .B2(_03604_),
    .ZN(_00374_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11451_ (.A1(\channels.accum[1][11] ),
    .A2(_03605_),
    .ZN(_03608_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11452_ (.A1(_03600_),
    .A2(_01459_),
    .B(_03608_),
    .ZN(_00375_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11453_ (.I(\channels.accum[1][12] ),
    .ZN(_03609_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11454_ (.A1(_03609_),
    .A2(_03603_),
    .B1(_01475_),
    .B2(_03604_),
    .ZN(_00376_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11455_ (.A1(\channels.accum[1][13] ),
    .A2(_03605_),
    .ZN(_03610_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11456_ (.A1(_03600_),
    .A2(_01487_),
    .B(_03610_),
    .ZN(_00377_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11457_ (.I(\channels.accum[1][14] ),
    .ZN(_03611_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11458_ (.A1(_03611_),
    .A2(_03603_),
    .B1(_01503_),
    .B2(_03604_),
    .ZN(_00378_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11459_ (.I(_02364_),
    .Z(_03612_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11460_ (.A1(\channels.accum[1][15] ),
    .A2(_03605_),
    .ZN(_03613_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11461_ (.A1(_03612_),
    .A2(_01515_),
    .B(_03613_),
    .ZN(_00379_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11462_ (.I(\channels.accum[1][16] ),
    .ZN(_03614_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11463_ (.I(_01104_),
    .Z(_03615_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11464_ (.I(_01219_),
    .Z(_03616_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11465_ (.A1(_03614_),
    .A2(_03615_),
    .B1(_01524_),
    .B2(_03616_),
    .ZN(_00380_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11466_ (.A1(\channels.accum[1][17] ),
    .A2(_01230_),
    .B1(_01530_),
    .B2(_01101_),
    .ZN(_03617_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11467_ (.I(_03617_),
    .ZN(_00381_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11468_ (.I(\channels.accum[1][18] ),
    .ZN(_03618_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11469_ (.A1(_03618_),
    .A2(_03615_),
    .B1(_01539_),
    .B2(_03616_),
    .ZN(_00382_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11470_ (.A1(\channels.accum[1][19] ),
    .A2(_03590_),
    .ZN(_03619_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11471_ (.A1(_03612_),
    .A2(_01545_),
    .B(_03619_),
    .ZN(_00383_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11472_ (.I(\channels.accum[1][20] ),
    .ZN(_03620_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11473_ (.A1(_03620_),
    .A2(_03615_),
    .B1(_01552_),
    .B2(_03616_),
    .ZN(_00384_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11474_ (.A1(\channels.accum[1][21] ),
    .A2(_03590_),
    .ZN(_03621_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11475_ (.A1(_03612_),
    .A2(_01559_),
    .B(_03621_),
    .ZN(_00385_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11476_ (.A1(_01563_),
    .A2(_03615_),
    .B1(_01568_),
    .B2(_03616_),
    .ZN(_00386_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11477_ (.A1(\channels.accum[1][23] ),
    .A2(_03590_),
    .ZN(_03622_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11478_ (.A1(_03612_),
    .A2(_01571_),
    .B(_03622_),
    .ZN(_00387_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11479_ (.A1(_00131_),
    .A2(_01033_),
    .B(_01029_),
    .ZN(_03623_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11480_ (.I(_03623_),
    .Z(_00389_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11481_ (.I(_00389_),
    .ZN(_00388_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11482_ (.A1(_02289_),
    .A2(_01954_),
    .Z(_03624_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11483_ (.I(_03624_),
    .Z(_03625_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11484_ (.I(_03624_),
    .Z(_03626_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11485_ (.I(_03516_),
    .Z(_03627_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11486_ (.A1(\channels.freq1[0] ),
    .A2(_03626_),
    .B(_03627_),
    .ZN(_03628_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11487_ (.A1(_02308_),
    .A2(_03625_),
    .B(_03628_),
    .ZN(_00390_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11488_ (.A1(\channels.freq1[1] ),
    .A2(_03626_),
    .B(_03627_),
    .ZN(_03629_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11489_ (.A1(_03511_),
    .A2(_03625_),
    .B(_03629_),
    .ZN(_00391_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11490_ (.A1(\channels.freq1[2] ),
    .A2(_03626_),
    .B(_03627_),
    .ZN(_03630_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11491_ (.A1(_03513_),
    .A2(_03625_),
    .B(_03630_),
    .ZN(_00392_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11492_ (.A1(\channels.freq1[3] ),
    .A2(_03626_),
    .B(_03627_),
    .ZN(_03631_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11493_ (.A1(_03515_),
    .A2(_03625_),
    .B(_03631_),
    .ZN(_00393_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11494_ (.I(_03624_),
    .Z(_03632_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11495_ (.I(_03624_),
    .Z(_03633_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11496_ (.I(_03516_),
    .Z(_03634_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11497_ (.A1(\channels.freq1[4] ),
    .A2(_03633_),
    .B(_03634_),
    .ZN(_03635_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11498_ (.A1(_02319_),
    .A2(_03632_),
    .B(_03635_),
    .ZN(_00394_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11499_ (.A1(\channels.freq1[5] ),
    .A2(_03633_),
    .B(_03634_),
    .ZN(_03636_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11500_ (.A1(_02324_),
    .A2(_03632_),
    .B(_03636_),
    .ZN(_00395_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11501_ (.A1(\channels.freq1[6] ),
    .A2(_03633_),
    .B(_03634_),
    .ZN(_03637_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11502_ (.A1(_02326_),
    .A2(_03632_),
    .B(_03637_),
    .ZN(_00396_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11503_ (.A1(\channels.freq1[7] ),
    .A2(_03633_),
    .B(_03634_),
    .ZN(_03638_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11504_ (.A1(_02328_),
    .A2(_03632_),
    .B(_03638_),
    .ZN(_00397_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11505_ (.I(_01740_),
    .Z(_03639_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11506_ (.I(_01779_),
    .Z(_03640_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11507_ (.A1(_03640_),
    .A2(_01885_),
    .Z(_03641_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11508_ (.I(_03641_),
    .Z(_03642_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11509_ (.I(_03641_),
    .Z(_03643_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11510_ (.I(_03516_),
    .Z(_03644_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11511_ (.A1(\channels.pw1[0] ),
    .A2(_03643_),
    .B(_03644_),
    .ZN(_03645_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11512_ (.A1(_03639_),
    .A2(_03642_),
    .B(_03645_),
    .ZN(_00398_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11513_ (.A1(\channels.pw1[1] ),
    .A2(_03643_),
    .B(_03644_),
    .ZN(_03646_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11514_ (.A1(_03511_),
    .A2(_03642_),
    .B(_03646_),
    .ZN(_00399_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11515_ (.A1(\channels.pw1[2] ),
    .A2(_03643_),
    .B(_03644_),
    .ZN(_03647_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11516_ (.A1(_03513_),
    .A2(_03642_),
    .B(_03647_),
    .ZN(_00400_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11517_ (.A1(\channels.pw1[3] ),
    .A2(_03643_),
    .B(_03644_),
    .ZN(_03648_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11518_ (.A1(_03515_),
    .A2(_03642_),
    .B(_03648_),
    .ZN(_00401_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11519_ (.I(_03641_),
    .Z(_03649_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11520_ (.I(_03641_),
    .Z(_03650_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11521_ (.I(_02333_),
    .Z(_03651_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11522_ (.I(_03651_),
    .Z(_03652_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11523_ (.A1(\channels.pw1[4] ),
    .A2(_03650_),
    .B(_03652_),
    .ZN(_03653_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11524_ (.A1(_02319_),
    .A2(_03649_),
    .B(_03653_),
    .ZN(_00402_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11525_ (.A1(\channels.pw1[5] ),
    .A2(_03650_),
    .B(_03652_),
    .ZN(_03654_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11526_ (.A1(_02324_),
    .A2(_03649_),
    .B(_03654_),
    .ZN(_00403_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11527_ (.A1(\channels.pw1[6] ),
    .A2(_03650_),
    .B(_03652_),
    .ZN(_03655_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11528_ (.A1(_02326_),
    .A2(_03649_),
    .B(_03655_),
    .ZN(_00404_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11529_ (.A1(\channels.pw1[7] ),
    .A2(_03650_),
    .B(_03652_),
    .ZN(_03656_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11530_ (.A1(_02328_),
    .A2(_03649_),
    .B(_03656_),
    .ZN(_00405_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11531_ (.A1(_03640_),
    .A2(_01880_),
    .Z(_03657_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11532_ (.I(_03657_),
    .Z(_03658_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11533_ (.I(_03657_),
    .Z(_03659_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11534_ (.I(_03651_),
    .Z(_03660_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11535_ (.A1(\channels.freq2[0] ),
    .A2(_03659_),
    .B(_03660_),
    .ZN(_03661_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11536_ (.A1(_03639_),
    .A2(_03658_),
    .B(_03661_),
    .ZN(_00406_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11537_ (.I(_01755_),
    .Z(_03662_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11538_ (.A1(\channels.freq2[1] ),
    .A2(_03659_),
    .B(_03660_),
    .ZN(_03663_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11539_ (.A1(_03662_),
    .A2(_03658_),
    .B(_03663_),
    .ZN(_00407_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11540_ (.I(_01765_),
    .Z(_03664_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11541_ (.A1(\channels.freq2[2] ),
    .A2(_03659_),
    .B(_03660_),
    .ZN(_03665_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11542_ (.A1(_03664_),
    .A2(_03658_),
    .B(_03665_),
    .ZN(_00408_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11543_ (.I(_02298_),
    .Z(_03666_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11544_ (.A1(\channels.freq2[3] ),
    .A2(_03659_),
    .B(_03660_),
    .ZN(_03667_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11545_ (.A1(_03666_),
    .A2(_03658_),
    .B(_03667_),
    .ZN(_00409_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11546_ (.I(_02149_),
    .Z(_03668_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11547_ (.I(_03657_),
    .Z(_03669_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11548_ (.I(_03657_),
    .Z(_03670_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11549_ (.I(_03651_),
    .Z(_03671_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11550_ (.A1(\channels.freq2[4] ),
    .A2(_03670_),
    .B(_03671_),
    .ZN(_03672_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11551_ (.A1(_03668_),
    .A2(_03669_),
    .B(_03672_),
    .ZN(_00410_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11552_ (.I(_02154_),
    .Z(_03673_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11553_ (.A1(\channels.freq2[5] ),
    .A2(_03670_),
    .B(_03671_),
    .ZN(_03674_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11554_ (.A1(_03673_),
    .A2(_03669_),
    .B(_03674_),
    .ZN(_00411_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11555_ (.I(_01812_),
    .Z(_03675_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11556_ (.A1(\channels.freq2[6] ),
    .A2(_03670_),
    .B(_03671_),
    .ZN(_03676_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11557_ (.A1(_03675_),
    .A2(_03669_),
    .B(_03676_),
    .ZN(_00412_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11558_ (.I(_01817_),
    .Z(_03677_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11559_ (.A1(\channels.freq2[7] ),
    .A2(_03670_),
    .B(_03671_),
    .ZN(_03678_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11560_ (.A1(_03677_),
    .A2(_03669_),
    .B(_03678_),
    .ZN(_00413_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11561_ (.A1(_03640_),
    .A2(_01871_),
    .Z(_03679_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11562_ (.I(_03679_),
    .Z(_03680_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11563_ (.I(_03679_),
    .Z(_03681_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11564_ (.I(_03651_),
    .Z(_03682_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11565_ (.A1(\channels.freq3[0] ),
    .A2(_03681_),
    .B(_03682_),
    .ZN(_03683_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11566_ (.A1(_03639_),
    .A2(_03680_),
    .B(_03683_),
    .ZN(_00414_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11567_ (.A1(\channels.freq3[1] ),
    .A2(_03681_),
    .B(_03682_),
    .ZN(_03684_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11568_ (.A1(_03662_),
    .A2(_03680_),
    .B(_03684_),
    .ZN(_00415_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11569_ (.A1(\channels.freq3[2] ),
    .A2(_03681_),
    .B(_03682_),
    .ZN(_03685_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11570_ (.A1(_03664_),
    .A2(_03680_),
    .B(_03685_),
    .ZN(_00416_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11571_ (.A1(\channels.freq3[3] ),
    .A2(_03681_),
    .B(_03682_),
    .ZN(_03686_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11572_ (.A1(_03666_),
    .A2(_03680_),
    .B(_03686_),
    .ZN(_00417_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11573_ (.I(_03679_),
    .Z(_03687_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11574_ (.I(_03679_),
    .Z(_03688_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11575_ (.I(_02333_),
    .Z(_03689_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11576_ (.I(_03689_),
    .Z(_03690_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11577_ (.A1(\channels.freq3[4] ),
    .A2(_03688_),
    .B(_03690_),
    .ZN(_03691_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11578_ (.A1(_03668_),
    .A2(_03687_),
    .B(_03691_),
    .ZN(_00418_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11579_ (.A1(\channels.freq3[5] ),
    .A2(_03688_),
    .B(_03690_),
    .ZN(_03692_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11580_ (.A1(_03673_),
    .A2(_03687_),
    .B(_03692_),
    .ZN(_00419_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11581_ (.A1(\channels.freq3[6] ),
    .A2(_03688_),
    .B(_03690_),
    .ZN(_03693_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11582_ (.A1(_03675_),
    .A2(_03687_),
    .B(_03693_),
    .ZN(_00420_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11583_ (.A1(\channels.freq3[7] ),
    .A2(_03688_),
    .B(_03690_),
    .ZN(_03694_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11584_ (.A1(_03677_),
    .A2(_03687_),
    .B(_03694_),
    .ZN(_00421_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11585_ (.A1(_03640_),
    .A2(_01896_),
    .Z(_03695_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11586_ (.I(_03695_),
    .Z(_03696_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11587_ (.I(_03695_),
    .Z(_03697_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11588_ (.I(_03689_),
    .Z(_03698_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11589_ (.A1(\channels.pw3[0] ),
    .A2(_03697_),
    .B(_03698_),
    .ZN(_03699_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11590_ (.A1(_03639_),
    .A2(_03696_),
    .B(_03699_),
    .ZN(_00422_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11591_ (.A1(\channels.pw3[1] ),
    .A2(_03697_),
    .B(_03698_),
    .ZN(_03700_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11592_ (.A1(_03662_),
    .A2(_03696_),
    .B(_03700_),
    .ZN(_00423_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11593_ (.A1(\channels.pw3[2] ),
    .A2(_03697_),
    .B(_03698_),
    .ZN(_03701_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11594_ (.A1(_03664_),
    .A2(_03696_),
    .B(_03701_),
    .ZN(_00424_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11595_ (.A1(\channels.pw3[3] ),
    .A2(_03697_),
    .B(_03698_),
    .ZN(_03702_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11596_ (.A1(_03666_),
    .A2(_03696_),
    .B(_03702_),
    .ZN(_00425_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11597_ (.I(_03695_),
    .Z(_03703_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11598_ (.I(_03695_),
    .Z(_03704_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11599_ (.I(_03689_),
    .Z(_03705_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11600_ (.A1(\channels.pw3[4] ),
    .A2(_03704_),
    .B(_03705_),
    .ZN(_03706_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11601_ (.A1(_03668_),
    .A2(_03703_),
    .B(_03706_),
    .ZN(_00426_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11602_ (.A1(\channels.pw3[5] ),
    .A2(_03704_),
    .B(_03705_),
    .ZN(_03707_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11603_ (.A1(_03673_),
    .A2(_03703_),
    .B(_03707_),
    .ZN(_00427_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11604_ (.A1(\channels.pw3[6] ),
    .A2(_03704_),
    .B(_03705_),
    .ZN(_03708_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11605_ (.A1(_03675_),
    .A2(_03703_),
    .B(_03708_),
    .ZN(_00428_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11606_ (.A1(\channels.pw3[7] ),
    .A2(_03704_),
    .B(_03705_),
    .ZN(_03709_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11607_ (.A1(_03677_),
    .A2(_03703_),
    .B(_03709_),
    .ZN(_00429_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11608_ (.I(_01740_),
    .Z(_03710_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11609_ (.A1(_01780_),
    .A2(_01848_),
    .Z(_03711_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11610_ (.I(_03711_),
    .Z(_03712_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11611_ (.I(_03711_),
    .Z(_03713_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11612_ (.I(_03689_),
    .Z(_03714_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11613_ (.A1(\channels.pw2[0] ),
    .A2(_03713_),
    .B(_03714_),
    .ZN(_03715_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11614_ (.A1(_03710_),
    .A2(_03712_),
    .B(_03715_),
    .ZN(_00430_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11615_ (.A1(\channels.pw2[1] ),
    .A2(_03713_),
    .B(_03714_),
    .ZN(_03716_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11616_ (.A1(_03662_),
    .A2(_03712_),
    .B(_03716_),
    .ZN(_00431_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11617_ (.A1(\channels.pw2[2] ),
    .A2(_03713_),
    .B(_03714_),
    .ZN(_03717_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11618_ (.A1(_03664_),
    .A2(_03712_),
    .B(_03717_),
    .ZN(_00432_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11619_ (.A1(\channels.pw2[3] ),
    .A2(_03713_),
    .B(_03714_),
    .ZN(_03718_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11620_ (.A1(_03666_),
    .A2(_03712_),
    .B(_03718_),
    .ZN(_00433_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11621_ (.I(_03711_),
    .Z(_03719_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11622_ (.I(_03711_),
    .Z(_03720_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11623_ (.I(_02100_),
    .Z(_03721_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11624_ (.I(_03721_),
    .Z(_03722_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11625_ (.A1(\channels.pw2[4] ),
    .A2(_03720_),
    .B(_03722_),
    .ZN(_03723_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11626_ (.A1(_03668_),
    .A2(_03719_),
    .B(_03723_),
    .ZN(_00434_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11627_ (.A1(\channels.pw2[5] ),
    .A2(_03720_),
    .B(_03722_),
    .ZN(_03724_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11628_ (.A1(_03673_),
    .A2(_03719_),
    .B(_03724_),
    .ZN(_00435_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11629_ (.A1(\channels.pw2[6] ),
    .A2(_03720_),
    .B(_03722_),
    .ZN(_03725_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11630_ (.A1(_03675_),
    .A2(_03719_),
    .B(_03725_),
    .ZN(_00436_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11631_ (.A1(\channels.pw2[7] ),
    .A2(_03720_),
    .B(_03722_),
    .ZN(_03726_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11632_ (.A1(_03677_),
    .A2(_03719_),
    .B(_03726_),
    .ZN(_00437_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11633_ (.A1(_01092_),
    .A2(_01093_),
    .ZN(_03727_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _11634_ (.I(_03727_),
    .Z(_03728_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11635_ (.I(_01068_),
    .Z(_03729_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11636_ (.I(_03729_),
    .Z(_03730_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11637_ (.I(_03730_),
    .Z(_03731_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11638_ (.I(_03731_),
    .Z(_03732_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11639_ (.I(_01750_),
    .Z(_03733_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11640_ (.I(_03733_),
    .Z(_03734_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11641_ (.I(_03734_),
    .Z(_03735_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11642_ (.A1(\channels.clk_div[0] ),
    .A2(_03732_),
    .B(_03735_),
    .ZN(_03736_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11643_ (.A1(_03728_),
    .A2(_03736_),
    .ZN(_00438_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _11644_ (.I(_01264_),
    .Z(_03737_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11645_ (.A1(_03737_),
    .A2(_03728_),
    .ZN(_03738_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _11646_ (.A1(_03737_),
    .A2(_03727_),
    .ZN(_03739_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11647_ (.A1(_02272_),
    .A2(_03739_),
    .ZN(_03740_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11648_ (.A1(_03738_),
    .A2(_03740_),
    .ZN(_00439_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11649_ (.A1(_01583_),
    .A2(_03739_),
    .Z(_03741_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11650_ (.A1(_01933_),
    .A2(_03741_),
    .ZN(_00440_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11651_ (.I(_02839_),
    .Z(_03742_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11652_ (.I(_03742_),
    .Z(_03743_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11653_ (.I(_01319_),
    .Z(_03744_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11654_ (.I(_03131_),
    .Z(_03745_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11655_ (.I(_03039_),
    .Z(_03746_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11656_ (.I(_02721_),
    .Z(_03747_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11657_ (.I(_02687_),
    .Z(_03748_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11658_ (.A1(_03748_),
    .A2(_03742_),
    .ZN(_03749_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11659_ (.A1(_03747_),
    .A2(_03749_),
    .ZN(_03750_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11660_ (.A1(_03746_),
    .A2(_03750_),
    .ZN(_03751_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _11661_ (.A1(_03096_),
    .A2(_03540_),
    .Z(_03752_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11662_ (.I(_03752_),
    .ZN(_03753_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11663_ (.A1(_03535_),
    .A2(_03751_),
    .A3(_03753_),
    .ZN(_03754_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _11664_ (.A1(_03745_),
    .A2(_03754_),
    .ZN(_03755_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11665_ (.A1(_03530_),
    .A2(_03531_),
    .ZN(_03756_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11666_ (.I(_03756_),
    .Z(_03757_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11667_ (.A1(\channels.sus_rel1[5] ),
    .A2(_01294_),
    .Z(_03758_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _11668_ (.A1(\channels.sus_rel3[5] ),
    .A2(_01081_),
    .B1(_01281_),
    .B2(\channels.sus_rel2[5] ),
    .C(_03758_),
    .ZN(_03759_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11669_ (.A1(_03540_),
    .A2(_03759_),
    .ZN(_03760_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _11670_ (.A1(_03748_),
    .A2(_03759_),
    .B(_03760_),
    .ZN(_03761_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11671_ (.A1(\channels.sus_rel1[4] ),
    .A2(_01294_),
    .Z(_03762_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _11672_ (.A1(\channels.sus_rel3[4] ),
    .A2(_01081_),
    .B1(_01281_),
    .B2(\channels.sus_rel2[4] ),
    .C(_03762_),
    .ZN(_03763_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11673_ (.I0(_02711_),
    .I1(_03539_),
    .S(_03763_),
    .Z(_03764_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11674_ (.A1(\channels.sus_rel3[7] ),
    .A2(_01080_),
    .Z(_03765_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _11675_ (.A1(\channels.sus_rel2[7] ),
    .A2(_01281_),
    .B1(_01295_),
    .B2(\channels.sus_rel1[7] ),
    .C(_03765_),
    .ZN(_03766_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11676_ (.A1(_01168_),
    .A2(_02532_),
    .ZN(_03767_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _11677_ (.A1(_01168_),
    .A2(_02533_),
    .B(_03767_),
    .ZN(_03768_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11678_ (.A1(\channels.sus_rel3[6] ),
    .A2(_01081_),
    .ZN(_03769_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11679_ (.A1(\channels.sus_rel2[6] ),
    .A2(_01280_),
    .B1(_01294_),
    .B2(\channels.sus_rel1[6] ),
    .ZN(_03770_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _11680_ (.A1(_03769_),
    .A2(_03770_),
    .ZN(_03771_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _11681_ (.A1(_03768_),
    .A2(_03088_),
    .B1(_03771_),
    .B2(_03747_),
    .ZN(_03772_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _11682_ (.A1(_03539_),
    .A2(_02711_),
    .B1(_03131_),
    .B2(_03766_),
    .C(_03772_),
    .ZN(_03773_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11683_ (.A1(_03748_),
    .A2(_02752_),
    .B1(_03766_),
    .B2(_03039_),
    .ZN(_03774_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11684_ (.A1(_03536_),
    .A2(_03535_),
    .ZN(_03775_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _11685_ (.A1(_03535_),
    .A2(_03771_),
    .B(_03774_),
    .C(_03775_),
    .ZN(_03776_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _11686_ (.A1(_03761_),
    .A2(_03764_),
    .A3(_03773_),
    .A4(_03776_),
    .ZN(_03777_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _11687_ (.A1(_03550_),
    .A2(_03755_),
    .B1(_03757_),
    .B2(_03777_),
    .ZN(_03778_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _11688_ (.A1(_03534_),
    .A2(_03778_),
    .Z(_03779_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11689_ (.I(_01425_),
    .Z(_03780_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11690_ (.A1(\channels.sus_rel3[0] ),
    .A2(_01439_),
    .B1(_03780_),
    .B2(\channels.sus_rel2[0] ),
    .ZN(_03781_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11691_ (.I(_01397_),
    .Z(_03782_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11692_ (.I(_01277_),
    .Z(_03783_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11693_ (.I(_03756_),
    .Z(_03784_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11694_ (.I(_03784_),
    .Z(_03785_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _11695_ (.A1(\channels.atk_dec3[0] ),
    .A2(_03782_),
    .B1(_03783_),
    .B2(\channels.atk_dec2[0] ),
    .C(_03785_),
    .ZN(_03786_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11696_ (.A1(_03757_),
    .A2(_03781_),
    .B(_03786_),
    .ZN(_03787_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11697_ (.I(_01290_),
    .Z(_03788_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11698_ (.I0(\channels.atk_dec1[0] ),
    .I1(\channels.sus_rel1[0] ),
    .S(_03784_),
    .Z(_03789_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11699_ (.A1(_03788_),
    .A2(_03789_),
    .Z(_03790_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11700_ (.I(_03532_),
    .Z(_03791_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _11701_ (.A1(\channels.atk_dec3[4] ),
    .A2(_01078_),
    .B1(_03780_),
    .B2(\channels.atk_dec2[4] ),
    .C1(_01291_),
    .C2(\channels.atk_dec1[4] ),
    .ZN(_03792_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11702_ (.A1(_03791_),
    .A2(_03792_),
    .ZN(_03793_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _11703_ (.A1(_03533_),
    .A2(_03787_),
    .A3(_03790_),
    .B(_03793_),
    .ZN(_03794_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11704_ (.A1(\channels.atk_dec3[1] ),
    .A2(_01077_),
    .B1(_01425_),
    .B2(\channels.atk_dec2[1] ),
    .ZN(_03795_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11705_ (.A1(\channels.sus_rel3[1] ),
    .A2(_01077_),
    .B1(_01425_),
    .B2(\channels.sus_rel2[1] ),
    .ZN(_03796_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11706_ (.I0(_03795_),
    .I1(_03796_),
    .S(_03785_),
    .Z(_03797_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11707_ (.I0(\channels.atk_dec1[1] ),
    .I1(\channels.sus_rel1[1] ),
    .S(_03784_),
    .Z(_03798_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11708_ (.A1(_03788_),
    .A2(_03798_),
    .B(_03532_),
    .ZN(_03799_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _11709_ (.A1(\channels.atk_dec3[5] ),
    .A2(_01078_),
    .B1(_03780_),
    .B2(\channels.atk_dec2[5] ),
    .C1(_01291_),
    .C2(\channels.atk_dec1[5] ),
    .ZN(_03800_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _11710_ (.A1(_03797_),
    .A2(_03799_),
    .B1(_03800_),
    .B2(_03791_),
    .ZN(_03801_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11711_ (.I(_03801_),
    .ZN(_03802_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11712_ (.I(_03802_),
    .Z(_03803_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _11713_ (.A1(_03794_),
    .A2(_03803_),
    .ZN(_03804_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11714_ (.I(_03794_),
    .ZN(_03805_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11715_ (.A1(\channels.sus_rel3[2] ),
    .A2(_03782_),
    .B1(_01278_),
    .B2(\channels.sus_rel2[2] ),
    .ZN(_03806_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _11716_ (.A1(\channels.atk_dec3[2] ),
    .A2(_03782_),
    .B1(_01278_),
    .B2(\channels.atk_dec2[2] ),
    .C(_03785_),
    .ZN(_03807_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _11717_ (.A1(_03757_),
    .A2(_03806_),
    .B(_03807_),
    .ZN(_03808_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11718_ (.I0(\channels.atk_dec1[2] ),
    .I1(\channels.sus_rel1[2] ),
    .S(_03784_),
    .Z(_03809_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11719_ (.A1(_03788_),
    .A2(_03809_),
    .Z(_03810_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _11720_ (.A1(\channels.atk_dec3[6] ),
    .A2(_01439_),
    .B1(_03783_),
    .B2(\channels.atk_dec2[6] ),
    .C1(_01291_),
    .C2(\channels.atk_dec1[6] ),
    .ZN(_03811_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11721_ (.A1(_03791_),
    .A2(_03811_),
    .ZN(_03812_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _11722_ (.A1(_03533_),
    .A2(_03808_),
    .A3(_03810_),
    .B(_03812_),
    .ZN(_03813_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _11723_ (.I(_03813_),
    .ZN(_03814_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11724_ (.A1(_03805_),
    .A2(_03814_),
    .ZN(_03815_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11725_ (.A1(_03803_),
    .A2(_03815_),
    .ZN(_03816_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11726_ (.A1(\channels.atk_dec3[3] ),
    .A2(_01439_),
    .B1(_03783_),
    .B2(\channels.atk_dec2[3] ),
    .ZN(_03817_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11727_ (.A1(\channels.sus_rel3[3] ),
    .A2(_03782_),
    .B1(_03783_),
    .B2(\channels.sus_rel2[3] ),
    .ZN(_03818_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11728_ (.I0(_03817_),
    .I1(_03818_),
    .S(_03757_),
    .Z(_03819_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11729_ (.I0(\channels.atk_dec1[3] ),
    .I1(\channels.sus_rel1[3] ),
    .S(_03785_),
    .Z(_03820_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11730_ (.A1(_01292_),
    .A2(_03820_),
    .B(_03791_),
    .ZN(_03821_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _11731_ (.A1(\channels.atk_dec3[7] ),
    .A2(_01078_),
    .B1(_03780_),
    .B2(\channels.atk_dec2[7] ),
    .C1(_03788_),
    .C2(\channels.atk_dec1[7] ),
    .ZN(_03822_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _11732_ (.A1(_03819_),
    .A2(_03821_),
    .B1(_03822_),
    .B2(_03533_),
    .ZN(_03823_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11733_ (.I(_03823_),
    .ZN(_03824_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11734_ (.A1(_03814_),
    .A2(_03824_),
    .ZN(_03825_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11735_ (.A1(_03813_),
    .A2(_03823_),
    .ZN(_03826_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11736_ (.A1(_03825_),
    .A2(_03826_),
    .ZN(_03827_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11737_ (.A1(_03801_),
    .A2(_03814_),
    .ZN(_03828_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11738_ (.A1(_03816_),
    .A2(_03827_),
    .B(_03828_),
    .ZN(_03829_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _11739_ (.A1(_03804_),
    .A2(_03829_),
    .ZN(_03830_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11740_ (.I(_01150_),
    .Z(_03831_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _11741_ (.I(_03831_),
    .Z(_03832_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _11742_ (.I0(\channels.env_counter[0][2] ),
    .I1(\channels.env_counter[1][2] ),
    .I2(\channels.env_counter[2][2] ),
    .I3(\channels.env_counter[3][2] ),
    .S0(_03832_),
    .S1(_01171_),
    .Z(_03833_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _11743_ (.A1(_03830_),
    .A2(_03833_),
    .Z(_03834_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11744_ (.I(_03823_),
    .Z(_03835_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11745_ (.I(_03835_),
    .Z(_03836_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11746_ (.I(_03794_),
    .Z(_03837_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11747_ (.A1(_03802_),
    .A2(_03813_),
    .ZN(_03838_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11748_ (.A1(_03828_),
    .A2(_03838_),
    .ZN(_03839_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11749_ (.A1(_03837_),
    .A2(_03839_),
    .Z(_03840_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11750_ (.A1(_03836_),
    .A2(_03840_),
    .ZN(_03841_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11751_ (.I(_01166_),
    .Z(_03842_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _11752_ (.I0(\channels.env_counter[0][9] ),
    .I1(\channels.env_counter[1][9] ),
    .I2(\channels.env_counter[2][9] ),
    .I3(\channels.env_counter[3][9] ),
    .S0(_03832_),
    .S1(_03842_),
    .Z(_03843_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11753_ (.A1(_03841_),
    .A2(_03843_),
    .Z(_03844_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11754_ (.I(_03813_),
    .Z(_03845_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11755_ (.A1(_03845_),
    .A2(_03835_),
    .ZN(_03846_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11756_ (.A1(_03805_),
    .A2(_03835_),
    .ZN(_03847_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11757_ (.A1(_03846_),
    .A2(_03847_),
    .ZN(_03848_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11758_ (.I(_03848_),
    .ZN(_03849_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11759_ (.I(_03801_),
    .Z(_03850_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11760_ (.A1(_03837_),
    .A2(_03850_),
    .ZN(_03851_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11761_ (.A1(_03837_),
    .A2(_03839_),
    .B(_03824_),
    .ZN(_03852_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11762_ (.A1(_03849_),
    .A2(_03851_),
    .B(_03852_),
    .ZN(_03853_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _11763_ (.I0(\channels.env_counter[0][6] ),
    .I1(\channels.env_counter[1][6] ),
    .I2(\channels.env_counter[2][6] ),
    .I3(\channels.env_counter[3][6] ),
    .S0(_03832_),
    .S1(_03842_),
    .Z(_03854_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11764_ (.A1(_03853_),
    .A2(_03854_),
    .Z(_03855_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _11765_ (.A1(_03834_),
    .A2(_03844_),
    .A3(_03855_),
    .ZN(_03856_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11766_ (.I(_03815_),
    .Z(_03857_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11767_ (.I(_03857_),
    .ZN(_03858_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11768_ (.A1(_03837_),
    .A2(_03827_),
    .B(_03858_),
    .ZN(_03859_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _11769_ (.A1(_03850_),
    .A2(_03859_),
    .ZN(_03860_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _11770_ (.I0(\channels.env_counter[0][5] ),
    .I1(\channels.env_counter[1][5] ),
    .I2(\channels.env_counter[2][5] ),
    .I3(\channels.env_counter[3][5] ),
    .S0(_01152_),
    .S1(_01171_),
    .Z(_03861_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11771_ (.I(_03861_),
    .Z(_03862_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11772_ (.A1(_03860_),
    .A2(_03862_),
    .ZN(_03863_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11773_ (.A1(_03850_),
    .A2(_03845_),
    .B(_03805_),
    .ZN(_03864_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11774_ (.A1(_03836_),
    .A2(_03839_),
    .B(_03864_),
    .ZN(_03865_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _11775_ (.I0(\channels.env_counter[0][4] ),
    .I1(\channels.env_counter[1][4] ),
    .I2(\channels.env_counter[2][4] ),
    .I3(\channels.env_counter[3][4] ),
    .S0(_03831_),
    .S1(_01167_),
    .Z(_03866_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _11776_ (.A1(_03865_),
    .A2(_03866_),
    .ZN(_03867_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11777_ (.A1(_03794_),
    .A2(_03845_),
    .ZN(_03868_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11778_ (.A1(_03801_),
    .A2(_03868_),
    .ZN(_03869_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11779_ (.A1(_03804_),
    .A2(_03869_),
    .ZN(_03870_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11780_ (.A1(_03824_),
    .A2(_03870_),
    .ZN(_03871_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11781_ (.A1(_03804_),
    .A2(_03825_),
    .ZN(_03872_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11782_ (.A1(_03871_),
    .A2(_03872_),
    .ZN(_03873_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _11783_ (.I0(\channels.env_counter[0][1] ),
    .I1(\channels.env_counter[1][1] ),
    .I2(\channels.env_counter[2][1] ),
    .I3(\channels.env_counter[3][1] ),
    .S0(_03831_),
    .S1(_01167_),
    .Z(_03874_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11784_ (.A1(_03873_),
    .A2(_03874_),
    .ZN(_03875_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _11785_ (.A1(_03863_),
    .A2(_03867_),
    .A3(_03875_),
    .ZN(_03876_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11786_ (.A1(_03803_),
    .A2(_03858_),
    .B(_03868_),
    .ZN(_03877_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _11787_ (.A1(_03846_),
    .A2(_03851_),
    .B1(_03877_),
    .B2(_03836_),
    .ZN(_03878_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _11788_ (.I0(\channels.env_counter[0][0] ),
    .I1(\channels.env_counter[1][0] ),
    .I2(\channels.env_counter[2][0] ),
    .I3(\channels.env_counter[3][0] ),
    .S0(_01151_),
    .S1(_01167_),
    .Z(_03879_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11789_ (.I(_03879_),
    .Z(_03880_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11790_ (.A1(_03878_),
    .A2(_03880_),
    .Z(_03881_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11791_ (.A1(_03878_),
    .A2(_03880_),
    .ZN(_03882_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11792_ (.A1(_03873_),
    .A2(_03874_),
    .ZN(_03883_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11793_ (.I(_03848_),
    .Z(_03884_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11794_ (.A1(_03804_),
    .A2(_03845_),
    .ZN(_03885_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _11795_ (.I(_01149_),
    .Z(_03886_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _11796_ (.I0(\channels.env_counter[0][3] ),
    .I1(\channels.env_counter[1][3] ),
    .I2(\channels.env_counter[2][3] ),
    .I3(\channels.env_counter[3][3] ),
    .S0(_03886_),
    .S1(_01166_),
    .Z(_03887_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11797_ (.I(_03887_),
    .Z(_03888_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11798_ (.A1(_03884_),
    .A2(_03885_),
    .B(_03888_),
    .ZN(_03889_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11799_ (.I(_03835_),
    .Z(_03890_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _11800_ (.A1(_03890_),
    .A2(_03869_),
    .A3(_03838_),
    .ZN(_03891_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _11801_ (.I0(\channels.env_counter[0][10] ),
    .I1(\channels.env_counter[1][10] ),
    .I2(\channels.env_counter[2][10] ),
    .I3(\channels.env_counter[3][10] ),
    .S0(_03886_),
    .S1(_01170_),
    .Z(_03892_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _11802_ (.A1(_03884_),
    .A2(_03885_),
    .A3(_03887_),
    .B1(_03891_),
    .B2(_03892_),
    .ZN(_03893_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11803_ (.I(_03893_),
    .ZN(_03894_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11804_ (.A1(_03860_),
    .A2(_03861_),
    .B(_03889_),
    .C(_03894_),
    .ZN(_03895_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _11805_ (.A1(_03881_),
    .A2(_03882_),
    .A3(_03883_),
    .A4(_03895_),
    .Z(_03896_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11806_ (.A1(_03890_),
    .A2(_03838_),
    .ZN(_03897_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _11807_ (.I0(\channels.env_counter[0][11] ),
    .I1(\channels.env_counter[1][11] ),
    .I2(\channels.env_counter[2][11] ),
    .I3(\channels.env_counter[3][11] ),
    .S0(_01150_),
    .S1(_01165_),
    .Z(_03898_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _11808_ (.A1(_03857_),
    .A2(_03897_),
    .A3(_03898_),
    .Z(_03899_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11809_ (.I(_03898_),
    .Z(_03900_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _11810_ (.A1(_03857_),
    .A2(_03897_),
    .B(_03900_),
    .ZN(_03901_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _11811_ (.A1(_03803_),
    .A2(_03857_),
    .B1(_03826_),
    .B2(_03884_),
    .ZN(_03902_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _11812_ (.I0(\channels.env_counter[0][7] ),
    .I1(\channels.env_counter[1][7] ),
    .I2(\channels.env_counter[2][7] ),
    .I3(\channels.env_counter[3][7] ),
    .S0(_01151_),
    .S1(_03842_),
    .Z(_03903_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11813_ (.A1(_03902_),
    .A2(_03903_),
    .ZN(_03904_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _11814_ (.I0(\channels.env_counter[0][8] ),
    .I1(\channels.env_counter[1][8] ),
    .I2(\channels.env_counter[2][8] ),
    .I3(\channels.env_counter[3][8] ),
    .S0(_03832_),
    .S1(_01171_),
    .Z(_03905_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11815_ (.I(_03828_),
    .Z(_03906_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11816_ (.I0(_03906_),
    .I1(_03816_),
    .S(_03836_),
    .Z(_03907_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _11817_ (.A1(_03905_),
    .A2(_03907_),
    .Z(_03908_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _11818_ (.I0(\channels.env_counter[0][12] ),
    .I1(\channels.env_counter[1][12] ),
    .I2(\channels.env_counter[2][12] ),
    .I3(\channels.env_counter[3][12] ),
    .S0(_01150_),
    .S1(_01166_),
    .Z(_03909_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11819_ (.A1(_03906_),
    .A2(_03847_),
    .B(_03909_),
    .ZN(_03910_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11820_ (.I(_03909_),
    .Z(_03911_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _11821_ (.A1(_03906_),
    .A2(_03847_),
    .A3(_03911_),
    .Z(_03912_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _11822_ (.A1(_03904_),
    .A2(_03908_),
    .A3(_03910_),
    .A4(_03912_),
    .Z(_03913_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11823_ (.I(_03905_),
    .Z(_03914_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11824_ (.A1(_03890_),
    .A2(_03868_),
    .Z(_03915_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11825_ (.I0(\channels.env_counter[0][13] ),
    .I1(\channels.env_counter[1][13] ),
    .S(_03886_),
    .Z(_03916_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11826_ (.I(\channels.env_counter[2][13] ),
    .ZN(_03917_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11827_ (.A1(_03831_),
    .A2(\channels.env_counter[3][13] ),
    .ZN(_03918_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _11828_ (.A1(_01151_),
    .A2(_03917_),
    .B(_03918_),
    .C(_01170_),
    .ZN(_03919_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _11829_ (.A1(_03842_),
    .A2(_03916_),
    .B(_03919_),
    .ZN(_03920_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11830_ (.A1(_03915_),
    .A2(_03920_),
    .ZN(_03921_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11831_ (.A1(_03891_),
    .A2(_03892_),
    .ZN(_03922_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11832_ (.A1(_03915_),
    .A2(_03920_),
    .ZN(_03923_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11833_ (.A1(_03850_),
    .A2(_03814_),
    .A3(_03890_),
    .ZN(_03924_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _11834_ (.I0(\channels.env_counter[0][14] ),
    .I1(\channels.env_counter[1][14] ),
    .I2(\channels.env_counter[2][14] ),
    .I3(\channels.env_counter[3][14] ),
    .S0(_03886_),
    .S1(_01170_),
    .Z(_03925_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11835_ (.A1(_03924_),
    .A2(_03925_),
    .Z(_03926_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11836_ (.A1(_03924_),
    .A2(_03925_),
    .ZN(_03927_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _11837_ (.A1(_03923_),
    .A2(_03926_),
    .A3(_03927_),
    .ZN(_03928_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _11838_ (.A1(_01584_),
    .A2(_03921_),
    .A3(_03922_),
    .A4(_03928_),
    .ZN(_03929_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _11839_ (.A1(_03902_),
    .A2(_03903_),
    .Z(_03930_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11840_ (.I(_03930_),
    .ZN(_03931_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _11841_ (.A1(_03914_),
    .A2(_03907_),
    .B(_03929_),
    .C(_03931_),
    .ZN(_03932_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _11842_ (.A1(_03899_),
    .A2(_03901_),
    .A3(_03913_),
    .A4(_03932_),
    .ZN(_03933_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _11843_ (.A1(_03856_),
    .A2(_03876_),
    .A3(_03896_),
    .A4(_03933_),
    .ZN(_03934_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11844_ (.I(_03934_),
    .Z(_03935_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11845_ (.A1(_03779_),
    .A2(_03935_),
    .Z(_03936_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11846_ (.I(_03936_),
    .Z(_03937_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11847_ (.A1(_03744_),
    .A2(_03937_),
    .ZN(_03938_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11848_ (.I(_03938_),
    .Z(_03939_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _11849_ (.I(_01087_),
    .Z(_03940_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11850_ (.A1(_03744_),
    .A2(_03937_),
    .B(_03940_),
    .ZN(_03941_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11851_ (.I(_03941_),
    .Z(_03942_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11852_ (.A1(\channels.env_vol[0][0] ),
    .A2(_03942_),
    .ZN(_03943_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11853_ (.A1(_03743_),
    .A2(_03939_),
    .B(_03943_),
    .ZN(_00441_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11854_ (.A1(_03537_),
    .A2(_03749_),
    .ZN(_03944_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11855_ (.A1(_03778_),
    .A2(_03934_),
    .ZN(_03945_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11856_ (.I(_03945_),
    .Z(_03946_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11857_ (.I(_03946_),
    .Z(_03947_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11858_ (.A1(_03944_),
    .A2(_03947_),
    .Z(_03948_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11859_ (.A1(\channels.env_vol[0][1] ),
    .A2(_03942_),
    .ZN(_03949_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11860_ (.A1(_03939_),
    .A2(_03948_),
    .B(_03949_),
    .ZN(_00442_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11861_ (.A1(_03748_),
    .A2(_03743_),
    .ZN(_03950_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11862_ (.I(_03945_),
    .Z(_03951_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11863_ (.A1(_03749_),
    .A2(_03946_),
    .ZN(_03952_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11864_ (.A1(_03950_),
    .A2(_03951_),
    .B(_03952_),
    .ZN(_03953_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11865_ (.A1(_03747_),
    .A2(_03953_),
    .Z(_03954_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11866_ (.A1(\channels.env_vol[0][2] ),
    .A2(_03942_),
    .ZN(_03955_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11867_ (.A1(_03939_),
    .A2(_03954_),
    .B(_03955_),
    .ZN(_00443_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11868_ (.A1(_03536_),
    .A2(_03951_),
    .ZN(_03956_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11869_ (.A1(_03950_),
    .A2(_03951_),
    .B1(_03956_),
    .B2(_03750_),
    .ZN(_03957_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11870_ (.A1(_03768_),
    .A2(_03957_),
    .Z(_03958_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11871_ (.A1(\channels.env_vol[0][3] ),
    .A2(_03942_),
    .ZN(_03959_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11872_ (.A1(_03939_),
    .A2(_03958_),
    .B(_03959_),
    .ZN(_00444_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11873_ (.I(_03938_),
    .Z(_03960_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11874_ (.I(_03751_),
    .Z(_03961_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11875_ (.A1(_03538_),
    .A2(_03951_),
    .ZN(_03962_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11876_ (.A1(_03961_),
    .A2(_03947_),
    .B(_03962_),
    .ZN(_03963_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11877_ (.A1(_03539_),
    .A2(_03963_),
    .Z(_03964_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11878_ (.I(_03941_),
    .Z(_03965_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11879_ (.A1(\channels.env_vol[0][4] ),
    .A2(_03965_),
    .ZN(_03966_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11880_ (.A1(_03960_),
    .A2(_03964_),
    .B(_03966_),
    .ZN(_00445_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11881_ (.A1(_03542_),
    .A2(_03752_),
    .ZN(_03967_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11882_ (.A1(_02752_),
    .A2(_03538_),
    .B(_03967_),
    .ZN(_03968_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11883_ (.I(_03961_),
    .ZN(_03969_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11884_ (.A1(_03540_),
    .A2(_03969_),
    .ZN(_03970_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _11885_ (.A1(_03541_),
    .A2(_03752_),
    .ZN(_03971_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11886_ (.A1(_03961_),
    .A2(_03971_),
    .ZN(_03972_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11887_ (.A1(_03970_),
    .A2(_03972_),
    .B(_03947_),
    .ZN(_03973_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _11888_ (.A1(_03947_),
    .A2(_03968_),
    .B(_03973_),
    .ZN(_03974_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11889_ (.A1(\channels.env_vol[0][5] ),
    .A2(_03965_),
    .ZN(_03975_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11890_ (.A1(_03960_),
    .A2(_03974_),
    .B(_03975_),
    .ZN(_00446_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11891_ (.A1(_03961_),
    .A2(_03753_),
    .ZN(_03976_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11892_ (.I0(_03976_),
    .I1(_03542_),
    .S(_03946_),
    .Z(_03977_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _11893_ (.A1(_03128_),
    .A2(_03977_),
    .Z(_03978_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11894_ (.A1(\channels.env_vol[0][6] ),
    .A2(_03965_),
    .ZN(_03979_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11895_ (.A1(_03960_),
    .A2(_03978_),
    .B(_03979_),
    .ZN(_00447_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11896_ (.I0(_03754_),
    .I1(_03543_),
    .S(_03946_),
    .Z(_03980_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11897_ (.A1(_03745_),
    .A2(_03980_),
    .Z(_03981_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11898_ (.A1(\channels.env_vol[0][7] ),
    .A2(_03965_),
    .ZN(_03982_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11899_ (.A1(_03960_),
    .A2(_03981_),
    .B(_03982_),
    .ZN(_00448_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11900_ (.A1(_03878_),
    .A2(_03879_),
    .ZN(_03983_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11901_ (.A1(_03923_),
    .A2(_03926_),
    .ZN(_03984_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11902_ (.A1(_03983_),
    .A2(_03921_),
    .A3(_03984_),
    .ZN(_03985_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _11903_ (.A1(_03905_),
    .A2(_03907_),
    .B(_03985_),
    .C(_03882_),
    .ZN(_03986_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _11904_ (.A1(_03930_),
    .A2(_03904_),
    .A3(_03908_),
    .A4(_03986_),
    .Z(_03987_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11905_ (.A1(_03860_),
    .A2(_03861_),
    .B(_03883_),
    .ZN(_03988_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11906_ (.A1(_03860_),
    .A2(_03862_),
    .B(_03988_),
    .ZN(_03989_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11907_ (.A1(_03844_),
    .A2(_03867_),
    .A3(_03875_),
    .ZN(_03990_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11908_ (.A1(_03891_),
    .A2(_03892_),
    .B(_03899_),
    .ZN(_03991_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11909_ (.I(_03991_),
    .ZN(_03992_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _11910_ (.A1(_03884_),
    .A2(_03885_),
    .A3(_03888_),
    .Z(_03993_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11911_ (.A1(_03901_),
    .A2(_03922_),
    .ZN(_03994_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11912_ (.A1(_01584_),
    .A2(_03910_),
    .ZN(_03995_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _11913_ (.A1(_03906_),
    .A2(_03847_),
    .A3(_03911_),
    .ZN(_03996_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _11914_ (.A1(_03994_),
    .A2(_03995_),
    .A3(_03996_),
    .A4(_03927_),
    .ZN(_03997_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _11915_ (.A1(_03992_),
    .A2(_03889_),
    .A3(_03993_),
    .A4(_03997_),
    .Z(_03998_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11916_ (.A1(_03855_),
    .A2(_03998_),
    .ZN(_03999_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _11917_ (.A1(_03989_),
    .A2(_03990_),
    .A3(_03999_),
    .ZN(_04000_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _11918_ (.A1(_03834_),
    .A2(_03987_),
    .A3(_04000_),
    .ZN(_04001_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _11919_ (.A1(_01185_),
    .A2(_01191_),
    .A3(_01198_),
    .A4(_01223_),
    .ZN(_04002_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11920_ (.A1(_03534_),
    .A2(_04002_),
    .B(_01585_),
    .ZN(_04003_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _11921_ (.A1(_04001_),
    .A2(_04003_),
    .ZN(_04004_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11922_ (.I(_04004_),
    .Z(_04005_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11923_ (.A1(_02356_),
    .A2(_04005_),
    .ZN(_04006_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11924_ (.I(_04006_),
    .Z(_04007_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11925_ (.I(_04007_),
    .Z(_04008_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11926_ (.I(_03935_),
    .Z(_04009_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _11927_ (.A1(_03880_),
    .A2(_04009_),
    .Z(_04010_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _11928_ (.A1(_01581_),
    .A2(_04005_),
    .B(_01102_),
    .ZN(_04011_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11929_ (.I(_04011_),
    .Z(_04012_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11930_ (.I(_04012_),
    .Z(_04013_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11931_ (.A1(\channels.env_counter[2][0] ),
    .A2(_04013_),
    .ZN(_04014_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11932_ (.A1(_04008_),
    .A2(_04010_),
    .B(_04014_),
    .ZN(_00449_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11933_ (.A1(_03879_),
    .A2(_03874_),
    .Z(_04015_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11934_ (.A1(_03880_),
    .A2(_03874_),
    .ZN(_04016_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _11935_ (.A1(_04009_),
    .A2(_04015_),
    .A3(_04016_),
    .Z(_04017_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11936_ (.A1(\channels.env_counter[2][1] ),
    .A2(_04013_),
    .ZN(_04018_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11937_ (.A1(_04008_),
    .A2(_04017_),
    .B(_04018_),
    .ZN(_00450_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11938_ (.I(_04001_),
    .Z(_04019_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11939_ (.A1(_03833_),
    .A2(_04015_),
    .Z(_04020_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11940_ (.A1(_04019_),
    .A2(_04020_),
    .ZN(_04021_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11941_ (.A1(\channels.env_counter[2][2] ),
    .A2(_04013_),
    .ZN(_04022_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11942_ (.A1(_04008_),
    .A2(_04021_),
    .B(_04022_),
    .ZN(_00451_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _11943_ (.A1(_03833_),
    .A2(_03888_),
    .A3(_04015_),
    .Z(_04023_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11944_ (.A1(_03833_),
    .A2(_04015_),
    .B(_03888_),
    .ZN(_04024_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _11945_ (.A1(_04009_),
    .A2(_04023_),
    .A3(_04024_),
    .Z(_04025_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11946_ (.A1(\channels.env_counter[2][3] ),
    .A2(_04013_),
    .ZN(_04026_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11947_ (.A1(_04008_),
    .A2(_04025_),
    .B(_04026_),
    .ZN(_00452_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11948_ (.I(_04006_),
    .Z(_04027_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11949_ (.A1(_03866_),
    .A2(_04023_),
    .Z(_04028_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11950_ (.A1(_04019_),
    .A2(_04028_),
    .ZN(_04029_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11951_ (.I(_04011_),
    .Z(_04030_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11952_ (.A1(\channels.env_counter[2][4] ),
    .A2(_04030_),
    .ZN(_04031_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11953_ (.A1(_04027_),
    .A2(_04029_),
    .B(_04031_),
    .ZN(_00453_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _11954_ (.A1(_03862_),
    .A2(_03866_),
    .A3(_04023_),
    .Z(_04032_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11955_ (.A1(_03866_),
    .A2(_04023_),
    .B(_03862_),
    .ZN(_04033_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _11956_ (.A1(_04009_),
    .A2(_04032_),
    .A3(_04033_),
    .Z(_04034_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11957_ (.A1(\channels.env_counter[2][5] ),
    .A2(_04030_),
    .ZN(_04035_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11958_ (.A1(_04027_),
    .A2(_04034_),
    .B(_04035_),
    .ZN(_00454_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11959_ (.A1(_03854_),
    .A2(_04032_),
    .Z(_04036_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11960_ (.A1(_04019_),
    .A2(_04036_),
    .ZN(_04037_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11961_ (.A1(\channels.env_counter[2][6] ),
    .A2(_04030_),
    .ZN(_04038_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11962_ (.A1(_04027_),
    .A2(_04037_),
    .B(_04038_),
    .ZN(_00455_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _11963_ (.A1(_03903_),
    .A2(_03854_),
    .A3(_04032_),
    .Z(_04039_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11964_ (.A1(_03854_),
    .A2(_04032_),
    .B(_03903_),
    .ZN(_04040_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _11965_ (.A1(_03935_),
    .A2(_04039_),
    .A3(_04040_),
    .Z(_04041_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11966_ (.A1(\channels.env_counter[2][7] ),
    .A2(_04030_),
    .ZN(_04042_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11967_ (.A1(_04027_),
    .A2(_04041_),
    .B(_04042_),
    .ZN(_00456_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11968_ (.I(_04006_),
    .Z(_04043_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11969_ (.I(_04001_),
    .Z(_04044_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11970_ (.A1(_03914_),
    .A2(_04039_),
    .ZN(_04045_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _11971_ (.A1(_03914_),
    .A2(_04039_),
    .Z(_04046_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _11972_ (.A1(_04044_),
    .A2(_04045_),
    .A3(_04046_),
    .ZN(_04047_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11973_ (.I(_04011_),
    .Z(_04048_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11974_ (.A1(\channels.env_counter[2][8] ),
    .A2(_04048_),
    .ZN(_04049_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11975_ (.A1(_04043_),
    .A2(_04047_),
    .B(_04049_),
    .ZN(_00457_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _11976_ (.A1(_03843_),
    .A2(_04045_),
    .ZN(_04050_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11977_ (.A1(_04019_),
    .A2(_04050_),
    .ZN(_04051_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11978_ (.A1(\channels.env_counter[2][9] ),
    .A2(_04048_),
    .ZN(_04052_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11979_ (.A1(_04043_),
    .A2(_04051_),
    .B(_04052_),
    .ZN(_00458_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11980_ (.I(_03892_),
    .ZN(_04053_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11981_ (.A1(_03914_),
    .A2(_03843_),
    .A3(_04039_),
    .ZN(_04054_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11982_ (.A1(_04053_),
    .A2(_04054_),
    .Z(_04055_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11983_ (.A1(_04044_),
    .A2(_04055_),
    .ZN(_04056_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11984_ (.A1(\channels.env_counter[2][10] ),
    .A2(_04048_),
    .ZN(_04057_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11985_ (.A1(_04043_),
    .A2(_04056_),
    .B(_04057_),
    .ZN(_00459_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11986_ (.A1(_04053_),
    .A2(_04054_),
    .ZN(_04058_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11987_ (.A1(_03900_),
    .A2(_04058_),
    .ZN(_04059_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _11988_ (.A1(_03900_),
    .A2(_04058_),
    .Z(_04060_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _11989_ (.A1(_04001_),
    .A2(_04059_),
    .A3(_04060_),
    .ZN(_04061_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11990_ (.A1(\channels.env_counter[2][11] ),
    .A2(_04048_),
    .ZN(_04062_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11991_ (.A1(_04043_),
    .A2(_04061_),
    .B(_04062_),
    .ZN(_00460_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _11992_ (.A1(_03911_),
    .A2(_04059_),
    .ZN(_04063_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11993_ (.A1(_04044_),
    .A2(_04063_),
    .ZN(_04064_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11994_ (.A1(\channels.env_counter[2][12] ),
    .A2(_04012_),
    .ZN(_04065_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11995_ (.A1(_04007_),
    .A2(_04064_),
    .B(_04065_),
    .ZN(_00461_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _11996_ (.A1(_03900_),
    .A2(_03911_),
    .A3(_04058_),
    .ZN(_04066_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11997_ (.A1(_03920_),
    .A2(_04066_),
    .Z(_04067_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11998_ (.A1(_04044_),
    .A2(_04067_),
    .ZN(_04068_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11999_ (.A1(\channels.env_counter[2][13] ),
    .A2(_04012_),
    .ZN(_04069_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12000_ (.A1(_04007_),
    .A2(_04068_),
    .B(_04069_),
    .ZN(_00462_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12001_ (.A1(_03920_),
    .A2(_04066_),
    .ZN(_04070_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _12002_ (.A1(_03925_),
    .A2(_04070_),
    .B(_03935_),
    .ZN(_04071_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _12003_ (.A1(_03925_),
    .A2(_04070_),
    .B(_04071_),
    .ZN(_04072_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12004_ (.A1(\channels.env_counter[2][14] ),
    .A2(_04012_),
    .ZN(_04073_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12005_ (.A1(_04007_),
    .A2(_04072_),
    .B(_04073_),
    .ZN(_00463_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _12006_ (.A1(_02363_),
    .A2(_04005_),
    .ZN(_04074_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12007_ (.I(_04074_),
    .Z(_04075_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12008_ (.I(_04075_),
    .Z(_04076_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _12009_ (.A1(_03737_),
    .A2(_04004_),
    .B(_01032_),
    .ZN(_04077_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12010_ (.I(_04077_),
    .Z(_04078_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12011_ (.I(_04078_),
    .Z(_04079_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12012_ (.A1(\channels.env_counter[1][0] ),
    .A2(_04079_),
    .ZN(_04080_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12013_ (.A1(_04010_),
    .A2(_04076_),
    .B(_04080_),
    .ZN(_00464_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12014_ (.A1(\channels.env_counter[1][1] ),
    .A2(_04079_),
    .ZN(_04081_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12015_ (.A1(_04017_),
    .A2(_04076_),
    .B(_04081_),
    .ZN(_00465_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12016_ (.A1(\channels.env_counter[1][2] ),
    .A2(_04079_),
    .ZN(_04082_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12017_ (.A1(_04021_),
    .A2(_04076_),
    .B(_04082_),
    .ZN(_00466_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12018_ (.A1(\channels.env_counter[1][3] ),
    .A2(_04079_),
    .ZN(_04083_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12019_ (.A1(_04025_),
    .A2(_04076_),
    .B(_04083_),
    .ZN(_00467_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12020_ (.I(_04074_),
    .Z(_04084_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12021_ (.I(_04077_),
    .Z(_04085_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12022_ (.A1(\channels.env_counter[1][4] ),
    .A2(_04085_),
    .ZN(_04086_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12023_ (.A1(_04029_),
    .A2(_04084_),
    .B(_04086_),
    .ZN(_00468_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12024_ (.A1(\channels.env_counter[1][5] ),
    .A2(_04085_),
    .ZN(_04087_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12025_ (.A1(_04034_),
    .A2(_04084_),
    .B(_04087_),
    .ZN(_00469_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12026_ (.A1(\channels.env_counter[1][6] ),
    .A2(_04085_),
    .ZN(_04088_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12027_ (.A1(_04037_),
    .A2(_04084_),
    .B(_04088_),
    .ZN(_00470_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12028_ (.A1(\channels.env_counter[1][7] ),
    .A2(_04085_),
    .ZN(_04089_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12029_ (.A1(_04041_),
    .A2(_04084_),
    .B(_04089_),
    .ZN(_00471_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12030_ (.I(_04074_),
    .Z(_04090_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12031_ (.I(_04077_),
    .Z(_04091_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12032_ (.A1(\channels.env_counter[1][8] ),
    .A2(_04091_),
    .ZN(_04092_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12033_ (.A1(_04047_),
    .A2(_04090_),
    .B(_04092_),
    .ZN(_00472_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12034_ (.A1(\channels.env_counter[1][9] ),
    .A2(_04091_),
    .ZN(_04093_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12035_ (.A1(_04051_),
    .A2(_04090_),
    .B(_04093_),
    .ZN(_00473_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12036_ (.A1(\channels.env_counter[1][10] ),
    .A2(_04091_),
    .ZN(_04094_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12037_ (.A1(_04056_),
    .A2(_04090_),
    .B(_04094_),
    .ZN(_00474_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12038_ (.A1(\channels.env_counter[1][11] ),
    .A2(_04091_),
    .ZN(_04095_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12039_ (.A1(_04061_),
    .A2(_04090_),
    .B(_04095_),
    .ZN(_00475_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12040_ (.A1(\channels.env_counter[1][12] ),
    .A2(_04078_),
    .ZN(_04096_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12041_ (.A1(_04064_),
    .A2(_04075_),
    .B(_04096_),
    .ZN(_00476_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12042_ (.A1(\channels.env_counter[1][13] ),
    .A2(_04078_),
    .ZN(_04097_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12043_ (.A1(_04068_),
    .A2(_04075_),
    .B(_04097_),
    .ZN(_00477_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12044_ (.A1(\channels.env_counter[1][14] ),
    .A2(_04078_),
    .ZN(_04098_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12045_ (.A1(_04072_),
    .A2(_04075_),
    .B(_04098_),
    .ZN(_00478_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12046_ (.I(\channels.adsr_state[3][0] ),
    .Z(_04099_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12047_ (.I(_04099_),
    .Z(_00479_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12048_ (.I(\channels.adsr_state[3][1] ),
    .Z(_04100_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12049_ (.I(_04100_),
    .Z(_00480_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _12050_ (.A1(\clk_ctr[0] ),
    .A2(_02354_),
    .A3(_03732_),
    .ZN(_00481_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12051_ (.I(_02353_),
    .Z(_04101_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12052_ (.A1(_01063_),
    .A2(\clk_ctr[1] ),
    .Z(_04102_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _12053_ (.A1(_04101_),
    .A2(_03732_),
    .A3(_04102_),
    .ZN(_00482_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _12054_ (.A1(_03744_),
    .A2(_04005_),
    .ZN(_04103_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12055_ (.I(_04103_),
    .Z(_04104_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12056_ (.I(_04104_),
    .Z(_04105_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _12057_ (.A1(_01319_),
    .A2(_04004_),
    .B(_01032_),
    .ZN(_04106_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12058_ (.I(_04106_),
    .Z(_04107_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12059_ (.I(_04107_),
    .Z(_04108_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12060_ (.A1(\channels.env_counter[0][0] ),
    .A2(_04108_),
    .ZN(_04109_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12061_ (.A1(_04010_),
    .A2(_04105_),
    .B(_04109_),
    .ZN(_00483_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12062_ (.A1(\channels.env_counter[0][1] ),
    .A2(_04108_),
    .ZN(_04110_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12063_ (.A1(_04017_),
    .A2(_04105_),
    .B(_04110_),
    .ZN(_00484_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12064_ (.A1(\channels.env_counter[0][2] ),
    .A2(_04108_),
    .ZN(_04111_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12065_ (.A1(_04021_),
    .A2(_04105_),
    .B(_04111_),
    .ZN(_00485_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12066_ (.A1(\channels.env_counter[0][3] ),
    .A2(_04108_),
    .ZN(_04112_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12067_ (.A1(_04025_),
    .A2(_04105_),
    .B(_04112_),
    .ZN(_00486_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12068_ (.I(_04103_),
    .Z(_04113_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12069_ (.I(_04106_),
    .Z(_04114_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12070_ (.A1(\channels.env_counter[0][4] ),
    .A2(_04114_),
    .ZN(_04115_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12071_ (.A1(_04029_),
    .A2(_04113_),
    .B(_04115_),
    .ZN(_00487_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12072_ (.A1(\channels.env_counter[0][5] ),
    .A2(_04114_),
    .ZN(_04116_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12073_ (.A1(_04034_),
    .A2(_04113_),
    .B(_04116_),
    .ZN(_00488_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12074_ (.A1(\channels.env_counter[0][6] ),
    .A2(_04114_),
    .ZN(_04117_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12075_ (.A1(_04037_),
    .A2(_04113_),
    .B(_04117_),
    .ZN(_00489_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12076_ (.A1(\channels.env_counter[0][7] ),
    .A2(_04114_),
    .ZN(_04118_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12077_ (.A1(_04041_),
    .A2(_04113_),
    .B(_04118_),
    .ZN(_00490_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12078_ (.I(_04103_),
    .Z(_04119_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12079_ (.I(_04106_),
    .Z(_04120_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12080_ (.A1(\channels.env_counter[0][8] ),
    .A2(_04120_),
    .ZN(_04121_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12081_ (.A1(_04047_),
    .A2(_04119_),
    .B(_04121_),
    .ZN(_00491_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12082_ (.A1(\channels.env_counter[0][9] ),
    .A2(_04120_),
    .ZN(_04122_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12083_ (.A1(_04051_),
    .A2(_04119_),
    .B(_04122_),
    .ZN(_00492_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12084_ (.A1(\channels.env_counter[0][10] ),
    .A2(_04120_),
    .ZN(_04123_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12085_ (.A1(_04056_),
    .A2(_04119_),
    .B(_04123_),
    .ZN(_00493_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12086_ (.A1(\channels.env_counter[0][11] ),
    .A2(_04120_),
    .ZN(_04124_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12087_ (.A1(_04061_),
    .A2(_04119_),
    .B(_04124_),
    .ZN(_00494_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12088_ (.A1(\channels.env_counter[0][12] ),
    .A2(_04107_),
    .ZN(_04125_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12089_ (.A1(_04064_),
    .A2(_04104_),
    .B(_04125_),
    .ZN(_00495_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12090_ (.A1(\channels.env_counter[0][13] ),
    .A2(_04107_),
    .ZN(_04126_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12091_ (.A1(_04068_),
    .A2(_04104_),
    .B(_04126_),
    .ZN(_00496_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12092_ (.A1(\channels.env_counter[0][14] ),
    .A2(_04107_),
    .ZN(_04127_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12093_ (.A1(_04072_),
    .A2(_04104_),
    .B(_04127_),
    .ZN(_00497_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _12094_ (.A1(_01240_),
    .A2(_03551_),
    .B(_01931_),
    .ZN(_04128_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12095_ (.I0(_03545_),
    .I1(\channels.adsr_state[2][0] ),
    .S(_04128_),
    .Z(_04129_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12096_ (.I(_04129_),
    .Z(_00498_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12097_ (.I0(_03554_),
    .I1(\channels.adsr_state[2][1] ),
    .S(_04128_),
    .Z(_04130_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12098_ (.I(_04130_),
    .Z(_00499_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _12099_ (.A1(_01219_),
    .A2(_03551_),
    .B(_01931_),
    .ZN(_04131_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12100_ (.I0(_03545_),
    .I1(\channels.adsr_state[1][0] ),
    .S(_04131_),
    .Z(_04132_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12101_ (.I(_04132_),
    .Z(_00500_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12102_ (.I0(_03554_),
    .I1(\channels.adsr_state[1][1] ),
    .S(_04131_),
    .Z(_04133_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12103_ (.I(_04133_),
    .Z(_00501_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12104_ (.I(\channels.accum[3][0] ),
    .Z(_04134_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12105_ (.I(_04134_),
    .Z(_00502_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12106_ (.I(\channels.accum[3][1] ),
    .Z(_04135_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12107_ (.I(_04135_),
    .Z(_00503_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12108_ (.I(\channels.accum[3][2] ),
    .Z(_04136_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12109_ (.I(_04136_),
    .Z(_00504_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12110_ (.I(\channels.accum[3][3] ),
    .Z(_04137_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12111_ (.I(_04137_),
    .Z(_00505_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12112_ (.I(\channels.accum[3][4] ),
    .Z(_04138_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12113_ (.I(_04138_),
    .Z(_00506_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12114_ (.I(\channels.accum[3][5] ),
    .Z(_04139_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12115_ (.I(_04139_),
    .Z(_00507_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12116_ (.I(\channels.accum[3][6] ),
    .Z(_04140_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12117_ (.I(_04140_),
    .Z(_00508_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12118_ (.I(\channels.accum[3][7] ),
    .Z(_04141_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12119_ (.I(_04141_),
    .Z(_00509_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12120_ (.I(\channels.accum[3][8] ),
    .Z(_04142_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12121_ (.I(_04142_),
    .Z(_00510_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12122_ (.I(\channels.accum[3][9] ),
    .Z(_04143_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12123_ (.I(_04143_),
    .Z(_00511_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12124_ (.I(\channels.accum[3][10] ),
    .Z(_04144_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12125_ (.I(_04144_),
    .Z(_00512_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12126_ (.I(\channels.accum[3][11] ),
    .Z(_04145_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12127_ (.I(_04145_),
    .Z(_00513_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12128_ (.I(\channels.accum[3][12] ),
    .Z(_04146_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12129_ (.I(_04146_),
    .Z(_00514_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12130_ (.I(\channels.accum[3][13] ),
    .Z(_04147_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12131_ (.I(_04147_),
    .Z(_00515_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12132_ (.I(\channels.accum[3][14] ),
    .Z(_04148_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12133_ (.I(_04148_),
    .Z(_00516_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12134_ (.I(\channels.accum[3][15] ),
    .Z(_04149_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12135_ (.I(_04149_),
    .Z(_00517_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12136_ (.I(\channels.accum[3][16] ),
    .Z(_04150_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12137_ (.I(_04150_),
    .Z(_00518_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12138_ (.I(\channels.accum[3][17] ),
    .Z(_04151_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12139_ (.I(_04151_),
    .Z(_00519_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12140_ (.I(\channels.accum[3][18] ),
    .Z(_04152_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12141_ (.I(_04152_),
    .Z(_00520_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12142_ (.I(\channels.accum[3][19] ),
    .Z(_04153_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12143_ (.I(_04153_),
    .Z(_00521_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12144_ (.I(\channels.accum[3][20] ),
    .Z(_04154_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12145_ (.I(_04154_),
    .Z(_00522_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12146_ (.I(\channels.accum[3][21] ),
    .Z(_04155_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12147_ (.I(_04155_),
    .Z(_00523_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12148_ (.I(\channels.accum[3][22] ),
    .Z(_04156_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12149_ (.I(_04156_),
    .Z(_00524_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12150_ (.I(\channels.accum[3][23] ),
    .Z(_04157_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12151_ (.I(_04157_),
    .Z(_00525_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12152_ (.I(_01093_),
    .Z(_04158_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _12153_ (.A1(_04158_),
    .A2(_03226_),
    .ZN(_04159_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12154_ (.I(_04159_),
    .Z(_04160_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12155_ (.I(_04160_),
    .Z(_04161_));
 gf180mcu_fd_sc_mcu7t5v0__or4_4 _12156_ (.A1(_03190_),
    .A2(_03312_),
    .A3(_03196_),
    .A4(\filters.high[5] ),
    .Z(_04162_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12157_ (.I(_04162_),
    .Z(_04163_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12158_ (.I(_04163_),
    .Z(_04164_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _12159_ (.A1(_03317_),
    .A2(_04164_),
    .ZN(_04165_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _12160_ (.A1(_03189_),
    .A2(_03181_),
    .A3(_03195_),
    .ZN(_04166_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12161_ (.I(_04166_),
    .Z(_04167_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12162_ (.I(_04167_),
    .Z(_04168_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12163_ (.I(_04168_),
    .Z(_04169_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _12164_ (.I(_04169_),
    .Z(_04170_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _12165_ (.A1(\filters.res_lut[3] ),
    .A2(_04170_),
    .ZN(_04171_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _12166_ (.A1(_04165_),
    .A2(_04171_),
    .ZN(_04172_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12167_ (.A1(\filters.res_lut[1] ),
    .A2(_04167_),
    .Z(_04173_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12168_ (.I(_04173_),
    .Z(_04174_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12169_ (.I(_04174_),
    .Z(_04175_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12170_ (.I(_04175_),
    .Z(_04176_));
 gf180mcu_fd_sc_mcu7t5v0__or4_2 _12171_ (.A1(_03311_),
    .A2(_03312_),
    .A3(_03313_),
    .A4(\filters.high[6] ),
    .Z(_04177_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _12172_ (.A1(_03331_),
    .A2(_04177_),
    .Z(_04178_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _12173_ (.I(_04178_),
    .Z(_04179_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12174_ (.I(_04179_),
    .Z(_04180_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12175_ (.I(_04180_),
    .Z(_04181_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12176_ (.I(_04181_),
    .Z(_04182_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12177_ (.A1(_04176_),
    .A2(_04182_),
    .ZN(_04183_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _12178_ (.A1(\filters.res_lut[0] ),
    .A2(_04167_),
    .Z(_04184_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12179_ (.I(_04184_),
    .Z(_04185_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12180_ (.I(_04185_),
    .Z(_04186_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12181_ (.I(_04186_),
    .Z(_04187_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _12182_ (.I(_03183_),
    .Z(_04188_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _12183_ (.I(_04188_),
    .Z(_04189_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _12184_ (.A1(_03239_),
    .A2(_03203_),
    .A3(_04189_),
    .A4(_03343_),
    .ZN(_04190_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12185_ (.I(_04190_),
    .Z(_04191_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12186_ (.I(_04191_),
    .Z(_04192_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _12187_ (.A1(_03350_),
    .A2(_04187_),
    .A3(_04192_),
    .ZN(_04193_));
 gf180mcu_fd_sc_mcu7t5v0__or4_4 _12188_ (.A1(_03189_),
    .A2(_03192_),
    .A3(_03195_),
    .A4(\filters.high[3] ),
    .Z(_04194_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _12189_ (.I(_04194_),
    .Z(_04195_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12190_ (.I(_04195_),
    .Z(_04196_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12191_ (.I(_04196_),
    .Z(_04197_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _12192_ (.A1(\filters.res_lut[4] ),
    .A2(_04168_),
    .Z(_04198_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12193_ (.I(_04198_),
    .Z(_04199_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _12194_ (.I(_04199_),
    .Z(_04200_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12195_ (.I(_04200_),
    .Z(_04201_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _12196_ (.A1(_03288_),
    .A2(_04197_),
    .A3(_04201_),
    .ZN(_04202_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12197_ (.A1(_04193_),
    .A2(_04202_),
    .Z(_04203_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _12198_ (.A1(_04193_),
    .A2(_04202_),
    .Z(_04204_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12199_ (.A1(_04183_),
    .A2(_04203_),
    .B(_04204_),
    .ZN(_04205_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12200_ (.I(_04182_),
    .Z(_04206_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12201_ (.A1(\filters.res_lut[2] ),
    .A2(_04169_),
    .Z(_04207_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12202_ (.I(_04207_),
    .Z(_04208_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12203_ (.A1(_04206_),
    .A2(_04208_),
    .ZN(_04209_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _12204_ (.A1(_04205_),
    .A2(_04209_),
    .ZN(_04210_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12205_ (.I(_04208_),
    .Z(_04211_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _12206_ (.A1(_04206_),
    .A2(_04205_),
    .A3(_04211_),
    .Z(_04212_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _12207_ (.A1(_04172_),
    .A2(_04210_),
    .B(_04212_),
    .ZN(_04213_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _12208_ (.I(\filters.high[0] ),
    .ZN(_04214_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _12209_ (.A1(_03239_),
    .A2(_03203_),
    .A3(_04189_),
    .A4(_04214_),
    .ZN(_04215_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12210_ (.I(_04215_),
    .Z(_04216_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _12211_ (.I(_04166_),
    .Z(_04217_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12212_ (.I0(\filters.cutoff_lut[6] ),
    .I1(\filters.res_lut[6] ),
    .S(_04217_),
    .Z(_04218_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12213_ (.I(_04218_),
    .Z(_04219_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12214_ (.I(_04219_),
    .Z(_04220_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12215_ (.I(_04220_),
    .Z(_04221_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12216_ (.I(_04221_),
    .Z(_04222_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _12217_ (.A1(_03200_),
    .A2(_04216_),
    .A3(_04222_),
    .ZN(_04223_));
 gf180mcu_fd_sc_mcu7t5v0__or4_2 _12218_ (.A1(_03311_),
    .A2(_03379_),
    .A3(_03313_),
    .A4(\filters.high[1] ),
    .Z(_04224_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12219_ (.I(_04224_),
    .Z(_04225_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12220_ (.I(_04225_),
    .Z(_04226_));
 gf180mcu_fd_sc_mcu7t5v0__and2_4 _12221_ (.A1(\filters.res_lut[5] ),
    .A2(_04167_),
    .Z(_04227_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12222_ (.I(_04227_),
    .Z(_04228_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _12223_ (.I(_04228_),
    .Z(_04229_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12224_ (.I(_04229_),
    .Z(_04230_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12225_ (.I(_04230_),
    .Z(_04231_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _12226_ (.A1(_03255_),
    .A2(_04226_),
    .A3(_04231_),
    .ZN(_04232_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _12227_ (.A1(_04223_),
    .A2(_04232_),
    .ZN(_04233_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _12228_ (.A1(_03255_),
    .A2(_04226_),
    .A3(_04221_),
    .ZN(_04234_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12229_ (.I0(\filters.cutoff_lut[7] ),
    .I1(\filters.res_lut[7] ),
    .S(_04217_),
    .Z(_04235_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12230_ (.I(_04235_),
    .Z(_04236_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12231_ (.I(_04236_),
    .Z(_04237_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12232_ (.I(_04237_),
    .Z(_04238_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _12233_ (.A1(_03200_),
    .A2(_04216_),
    .A3(_04238_),
    .ZN(_04239_));
 gf180mcu_fd_sc_mcu7t5v0__or4_4 _12234_ (.A1(_03246_),
    .A2(_03193_),
    .A3(_03249_),
    .A4(\filters.high[2] ),
    .Z(_04240_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _12235_ (.I(_04240_),
    .Z(_04241_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12236_ (.I(_04241_),
    .Z(_04242_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12237_ (.I(_04242_),
    .Z(_04243_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _12238_ (.A1(_03273_),
    .A2(_04243_),
    .A3(_04231_),
    .Z(_04244_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _12239_ (.A1(_04234_),
    .A2(_04239_),
    .A3(_04244_),
    .Z(_04245_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12240_ (.A1(_04233_),
    .A2(_04245_),
    .ZN(_04246_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _12241_ (.A1(_04183_),
    .A2(_04193_),
    .A3(_04202_),
    .Z(_04247_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12242_ (.A1(_04233_),
    .A2(_04245_),
    .ZN(_04248_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _12243_ (.A1(_04246_),
    .A2(_04247_),
    .B(_04248_),
    .ZN(_04249_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12244_ (.A1(_04234_),
    .A2(_04239_),
    .ZN(_04250_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12245_ (.A1(_04234_),
    .A2(_04239_),
    .ZN(_04251_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _12246_ (.A1(_04244_),
    .A2(_04250_),
    .B(_04251_),
    .ZN(_04252_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _12247_ (.I(_04235_),
    .Z(_04253_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _12248_ (.I(_04253_),
    .Z(_04254_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _12249_ (.I(_04254_),
    .Z(_04255_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _12250_ (.A1(_03254_),
    .A2(_04226_),
    .A3(_04255_),
    .ZN(_04256_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12251_ (.I(_04218_),
    .Z(_04257_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _12252_ (.I(_04257_),
    .Z(_04258_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _12253_ (.I(_04258_),
    .Z(_04259_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _12254_ (.A1(_03272_),
    .A2(_04243_),
    .A3(_04259_),
    .ZN(_04260_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _12255_ (.A1(_03288_),
    .A2(_04197_),
    .ZN(_04261_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12256_ (.A1(\filters.res_lut[5] ),
    .A2(_04168_),
    .ZN(_04262_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12257_ (.A1(_04261_),
    .A2(_04262_),
    .ZN(_04263_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _12258_ (.A1(_04256_),
    .A2(_04260_),
    .A3(_04263_),
    .ZN(_04264_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _12259_ (.I(_04174_),
    .Z(_04265_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12260_ (.I(_04265_),
    .Z(_04266_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _12261_ (.A1(_03348_),
    .A2(_04190_),
    .Z(_04267_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12262_ (.I(_04267_),
    .Z(_04268_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12263_ (.I(_04268_),
    .Z(_04269_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12264_ (.A1(_04266_),
    .A2(_04269_),
    .ZN(_04270_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _12265_ (.A1(_03238_),
    .A2(_03203_),
    .A3(_04188_),
    .A4(_03359_),
    .ZN(_04271_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _12266_ (.A1(_03362_),
    .A2(_04271_),
    .Z(_04272_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12267_ (.I(_04272_),
    .Z(_04273_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12268_ (.I(_04273_),
    .Z(_04274_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12269_ (.A1(_04274_),
    .A2(_04187_),
    .ZN(_04275_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _12270_ (.A1(_03180_),
    .A2(_03181_),
    .A3(_03183_),
    .A4(_03298_),
    .ZN(_04276_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12271_ (.A1(_03301_),
    .A2(_04276_),
    .Z(_04277_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12272_ (.I(_04277_),
    .Z(_04278_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12273_ (.I(_04278_),
    .Z(_04279_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12274_ (.I(_04279_),
    .Z(_04280_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12275_ (.I(_04280_),
    .Z(_04281_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12276_ (.A1(_04281_),
    .A2(_04201_),
    .ZN(_04282_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _12277_ (.A1(_04270_),
    .A2(_04275_),
    .A3(_04282_),
    .ZN(_04283_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _12278_ (.A1(_04252_),
    .A2(_04264_),
    .A3(_04283_),
    .Z(_04284_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12279_ (.A1(_04249_),
    .A2(_04284_),
    .ZN(_04285_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12280_ (.A1(\filters.res_lut[3] ),
    .A2(_04169_),
    .Z(_04286_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12281_ (.I(_04286_),
    .Z(_04287_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12282_ (.I(_04287_),
    .Z(_04288_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12283_ (.A1(_04206_),
    .A2(_04288_),
    .ZN(_04289_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12284_ (.I(_04273_),
    .Z(_04290_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12285_ (.I(_04290_),
    .Z(_04291_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12286_ (.I(_04291_),
    .Z(_04292_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12287_ (.I(_04187_),
    .Z(_04293_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12288_ (.I(_04198_),
    .Z(_04294_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12289_ (.I(_04294_),
    .Z(_04295_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12290_ (.I(_04295_),
    .Z(_04296_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12291_ (.I(_04281_),
    .Z(_04297_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _12292_ (.A1(_04292_),
    .A2(_04293_),
    .B1(_04296_),
    .B2(_04297_),
    .ZN(_04298_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _12293_ (.A1(_04281_),
    .A2(_04291_),
    .A3(_04293_),
    .A4(_04296_),
    .ZN(_04299_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12294_ (.A1(_04270_),
    .A2(_04298_),
    .B(_04299_),
    .ZN(_04300_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12295_ (.I(_04269_),
    .Z(_04301_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12296_ (.I(_04207_),
    .Z(_04302_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12297_ (.A1(_04301_),
    .A2(_04302_),
    .ZN(_04303_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12298_ (.A1(_04300_),
    .A2(_04303_),
    .Z(_04304_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12299_ (.A1(_04289_),
    .A2(_04304_),
    .Z(_04305_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12300_ (.A1(_04285_),
    .A2(_04305_),
    .Z(_04306_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _12301_ (.A1(_04249_),
    .A2(_04284_),
    .A3(_04305_),
    .ZN(_04307_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12302_ (.A1(_04213_),
    .A2(_04306_),
    .B(_04307_),
    .ZN(_04308_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _12303_ (.I(_04308_),
    .ZN(_04309_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _12304_ (.A1(_04213_),
    .A2(_04306_),
    .ZN(_04310_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12305_ (.A1(_03199_),
    .A2(_04216_),
    .Z(_04311_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12306_ (.I(_04311_),
    .Z(_04312_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12307_ (.I(_04312_),
    .Z(_04313_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12308_ (.I0(\filters.cutoff_lut[9] ),
    .I1(\filters.res_lut[9] ),
    .S(_04217_),
    .Z(_04314_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12309_ (.I(_04314_),
    .Z(_04315_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12310_ (.I(_04315_),
    .Z(_04316_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12311_ (.I(_04316_),
    .Z(_04317_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12312_ (.I(_04317_),
    .Z(_04318_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _12313_ (.A1(_04313_),
    .A2(_04318_),
    .ZN(_04319_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _12314_ (.A1(_03253_),
    .A2(_04224_),
    .Z(_04320_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12315_ (.I(_04320_),
    .Z(_04321_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12316_ (.I(_04321_),
    .Z(_04322_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12317_ (.I0(\filters.cutoff_lut[8] ),
    .I1(\filters.res_lut[8] ),
    .S(_04217_),
    .Z(_04323_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12318_ (.I(_04323_),
    .Z(_04324_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12319_ (.I(_04324_),
    .Z(_04325_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12320_ (.I(_04325_),
    .Z(_04326_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _12321_ (.A1(_04322_),
    .A2(_04326_),
    .ZN(_04327_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _12322_ (.A1(_04319_),
    .A2(_04327_),
    .ZN(_04328_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12323_ (.A1(_04256_),
    .A2(_04260_),
    .ZN(_04329_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12324_ (.A1(_04256_),
    .A2(_04260_),
    .ZN(_04330_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _12325_ (.A1(_04263_),
    .A2(_04329_),
    .B(_04330_),
    .ZN(_04331_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12326_ (.I(_04276_),
    .Z(_04332_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12327_ (.A1(_03302_),
    .A2(_04332_),
    .ZN(_04333_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12328_ (.A1(_04262_),
    .A2(_04333_),
    .ZN(_04334_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _12329_ (.A1(_03271_),
    .A2(_04253_),
    .A3(_04241_),
    .ZN(_04335_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _12330_ (.A1(_03287_),
    .A2(_04219_),
    .A3(_04196_),
    .ZN(_04336_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12331_ (.A1(_04335_),
    .A2(_04336_),
    .Z(_04337_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _12332_ (.A1(_04334_),
    .A2(_04337_),
    .ZN(_04338_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _12333_ (.A1(_04331_),
    .A2(_04338_),
    .Z(_04339_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12334_ (.A1(_04291_),
    .A2(_04266_),
    .ZN(_04340_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _12335_ (.A1(_03238_),
    .A2(_03182_),
    .A3(_04188_),
    .A4(_03373_),
    .ZN(_04341_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12336_ (.I(_04341_),
    .Z(_04342_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _12337_ (.A1(_03383_),
    .A2(_04342_),
    .A3(_04185_),
    .ZN(_04343_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _12338_ (.A1(_03316_),
    .A2(_04164_),
    .A3(_04199_),
    .ZN(_04344_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _12339_ (.A1(_04343_),
    .A2(_04344_),
    .ZN(_04345_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _12340_ (.A1(_04345_),
    .A2(_04340_),
    .ZN(_04346_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _12341_ (.I(_04346_),
    .ZN(_04347_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12342_ (.A1(_04339_),
    .A2(_04347_),
    .Z(_04348_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12343_ (.A1(_04252_),
    .A2(_04264_),
    .ZN(_04349_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12344_ (.A1(_04252_),
    .A2(_04264_),
    .ZN(_04350_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _12345_ (.A1(_04349_),
    .A2(_04283_),
    .B(_04350_),
    .ZN(_04351_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _12346_ (.A1(_04328_),
    .A2(_04348_),
    .A3(_04351_),
    .Z(_04352_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12347_ (.I(_04313_),
    .Z(_04353_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12348_ (.I(_04353_),
    .Z(_04354_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12349_ (.I(_04325_),
    .Z(_04355_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _12350_ (.A1(_04354_),
    .A2(_04355_),
    .ZN(_04356_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _12351_ (.A1(_04252_),
    .A2(_04264_),
    .A3(_04283_),
    .ZN(_04357_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12352_ (.A1(_04357_),
    .A2(_04249_),
    .Z(_04358_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _12353_ (.A1(_04356_),
    .A2(_04358_),
    .ZN(_04359_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12354_ (.A1(_04352_),
    .A2(_04359_),
    .ZN(_04360_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12355_ (.A1(_04352_),
    .A2(_04359_),
    .ZN(_04361_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _12356_ (.A1(_04310_),
    .A2(_04360_),
    .B(_04361_),
    .ZN(_04362_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12357_ (.A1(_04348_),
    .A2(_04351_),
    .Z(_04363_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12358_ (.A1(_04328_),
    .A2(_04363_),
    .ZN(_04364_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12359_ (.A1(_04319_),
    .A2(_04327_),
    .ZN(_04365_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12360_ (.I(_04323_),
    .Z(_04366_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12361_ (.I(_04366_),
    .Z(_04367_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _12362_ (.A1(_04241_),
    .A2(_03270_),
    .Z(_04368_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12363_ (.I(_04368_),
    .Z(_04369_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12364_ (.A1(_04367_),
    .A2(_04369_),
    .ZN(_04370_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12365_ (.I(_04314_),
    .Z(_04371_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12366_ (.I(_04371_),
    .Z(_04372_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12367_ (.A1(_04372_),
    .A2(_04321_),
    .ZN(_04373_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12368_ (.I0(\filters.cutoff_lut[10] ),
    .I1(\filters.res_lut[10] ),
    .S(_04166_),
    .Z(_04374_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12369_ (.I(_04374_),
    .Z(_04375_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12370_ (.I(_04375_),
    .Z(_04376_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12371_ (.I(_04376_),
    .Z(_04377_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12372_ (.I(_04377_),
    .Z(_04378_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12373_ (.A1(_04312_),
    .A2(_04378_),
    .ZN(_04379_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _12374_ (.A1(_04370_),
    .A2(_04373_),
    .A3(_04379_),
    .Z(_04380_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _12375_ (.A1(_04365_),
    .A2(_04380_),
    .Z(_04381_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12376_ (.A1(_04335_),
    .A2(_04336_),
    .ZN(_04382_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _12377_ (.A1(_04334_),
    .A2(_04337_),
    .B(_04382_),
    .ZN(_04383_));
 gf180mcu_fd_sc_mcu7t5v0__and2_4 _12378_ (.A1(_04162_),
    .A2(_03315_),
    .Z(_04384_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _12379_ (.I(_04384_),
    .Z(_04385_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _12380_ (.I(_04385_),
    .Z(_04386_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _12381_ (.A1(_04229_),
    .A2(_04386_),
    .ZN(_04387_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _12382_ (.I(_04253_),
    .Z(_04388_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _12383_ (.A1(_03286_),
    .A2(_04195_),
    .Z(_04389_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12384_ (.I(_04389_),
    .Z(_04390_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _12385_ (.A1(_04388_),
    .A2(_04390_),
    .ZN(_04391_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12386_ (.I(_04258_),
    .Z(_04392_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12387_ (.A1(_04392_),
    .A2(_04280_),
    .ZN(_04393_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _12388_ (.A1(_04387_),
    .A2(_04391_),
    .A3(_04393_),
    .Z(_04394_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _12389_ (.A1(_03381_),
    .A2(_04341_),
    .Z(_04395_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12390_ (.I(_04395_),
    .Z(_04396_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12391_ (.I(_04396_),
    .Z(_04397_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12392_ (.A1(_04265_),
    .A2(_04397_),
    .ZN(_04398_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12393_ (.A1(_04200_),
    .A2(_04181_),
    .ZN(_04399_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12394_ (.I(_04184_),
    .Z(_04400_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12395_ (.I(_04400_),
    .Z(_04401_));
 gf180mcu_fd_sc_mcu7t5v0__or4_2 _12396_ (.A1(_03190_),
    .A2(_03312_),
    .A3(_03196_),
    .A4(\filters.high[10] ),
    .Z(_04402_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _12397_ (.I(_04402_),
    .Z(_04403_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12398_ (.A1(_03398_),
    .A2(_04403_),
    .Z(_04404_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12399_ (.I(_04404_),
    .Z(_04405_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12400_ (.I(_04405_),
    .Z(_04406_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12401_ (.A1(_04401_),
    .A2(_04406_),
    .ZN(_04407_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _12402_ (.A1(_04398_),
    .A2(_04399_),
    .A3(_04407_),
    .Z(_04408_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _12403_ (.A1(_04383_),
    .A2(_04394_),
    .A3(_04408_),
    .ZN(_04409_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _12404_ (.I(_04409_),
    .ZN(_04410_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12405_ (.A1(_04331_),
    .A2(_04338_),
    .ZN(_04411_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _12406_ (.A1(_04339_),
    .A2(_04347_),
    .B(_04411_),
    .ZN(_04412_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _12407_ (.A1(_04381_),
    .A2(_04410_),
    .A3(_04412_),
    .Z(_04413_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12408_ (.A1(_04339_),
    .A2(net34),
    .Z(_04414_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _12409_ (.A1(_04414_),
    .A2(_04351_),
    .Z(_04415_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _12410_ (.I(_04302_),
    .Z(_04416_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _12411_ (.A1(_04301_),
    .A2(_04416_),
    .A3(_04300_),
    .Z(_04417_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12412_ (.A1(_04289_),
    .A2(_04304_),
    .ZN(_04418_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12413_ (.A1(_04417_),
    .A2(_04418_),
    .ZN(_04419_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12414_ (.I(_04287_),
    .Z(_04420_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12415_ (.A1(_04301_),
    .A2(_04420_),
    .ZN(_04421_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _12416_ (.A1(_04343_),
    .A2(_04344_),
    .Z(_04422_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12417_ (.A1(_04340_),
    .A2(_04345_),
    .B(_04422_),
    .ZN(_04423_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12418_ (.A1(_04292_),
    .A2(_04208_),
    .ZN(_04424_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _12419_ (.A1(_04423_),
    .A2(_04424_),
    .ZN(_04425_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _12420_ (.A1(_04421_),
    .A2(_04425_),
    .ZN(_04426_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _12421_ (.A1(_04415_),
    .A2(_04419_),
    .A3(_04426_),
    .Z(_04427_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _12422_ (.A1(_04364_),
    .A2(_04413_),
    .A3(_04427_),
    .ZN(_04428_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _12423_ (.A1(_04362_),
    .A2(_04428_),
    .ZN(_04429_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12424_ (.A1(_04362_),
    .A2(_04428_),
    .ZN(_04430_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _12425_ (.A1(_04309_),
    .A2(_04429_),
    .B(_04430_),
    .ZN(_04431_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _12426_ (.I(_04415_),
    .ZN(_04432_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12427_ (.A1(_04415_),
    .A2(_04426_),
    .Z(_04433_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12428_ (.A1(_04419_),
    .A2(_04433_),
    .ZN(_04434_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _12429_ (.A1(_04432_),
    .A2(_04426_),
    .B(_04434_),
    .ZN(_04435_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12430_ (.A1(_04328_),
    .A2(_04363_),
    .B(_04413_),
    .ZN(_04436_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _12431_ (.A1(_04328_),
    .A2(_04363_),
    .A3(_04413_),
    .ZN(_04437_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _12432_ (.A1(_04436_),
    .A2(_04427_),
    .B(_04437_),
    .ZN(_04438_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12433_ (.A1(net33),
    .A2(_04412_),
    .Z(_04439_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12434_ (.A1(_04381_),
    .A2(_04439_),
    .ZN(_04440_));
 gf180mcu_fd_sc_mcu7t5v0__or3_4 _12435_ (.A1(\filters.filter_step[2] ),
    .A2(_03181_),
    .A3(\filters.filter_step[0] ),
    .Z(_04441_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12436_ (.I(_04441_),
    .Z(_04442_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12437_ (.A1(\filters.cutoff_lut[11] ),
    .A2(_04442_),
    .Z(_04443_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12438_ (.I(_04443_),
    .Z(_04444_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12439_ (.I(_04444_),
    .Z(_04445_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12440_ (.I(_04445_),
    .Z(_04446_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12441_ (.I(_04446_),
    .Z(_04447_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _12442_ (.A1(_04353_),
    .A2(_04447_),
    .ZN(_04448_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12443_ (.I(_04372_),
    .Z(_04449_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _12444_ (.I(_04375_),
    .Z(_04450_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12445_ (.I(_04450_),
    .Z(_04451_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12446_ (.I(_04451_),
    .Z(_04452_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12447_ (.I(_04452_),
    .Z(_04453_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _12448_ (.A1(_04449_),
    .A2(_04322_),
    .B1(_04453_),
    .B2(_04312_),
    .ZN(_04454_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _12449_ (.A1(_04312_),
    .A2(_04449_),
    .A3(_04321_),
    .A4(_04453_),
    .ZN(_04455_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _12450_ (.A1(_04370_),
    .A2(_04454_),
    .B(_04455_),
    .ZN(_04456_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12451_ (.A1(_04366_),
    .A2(_04390_),
    .Z(_04457_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _12452_ (.A1(_03254_),
    .A2(_04225_),
    .A3(_04376_),
    .ZN(_04458_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _12453_ (.A1(_03273_),
    .A2(_04372_),
    .A3(_04243_),
    .ZN(_04459_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _12454_ (.A1(_04457_),
    .A2(_04458_),
    .A3(_04459_),
    .Z(_04460_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _12455_ (.A1(_04456_),
    .A2(_04460_),
    .ZN(_04461_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12456_ (.A1(_04448_),
    .A2(_04461_),
    .Z(_04462_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12457_ (.A1(_04383_),
    .A2(_04394_),
    .Z(_04463_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _12458_ (.A1(_04383_),
    .A2(_04394_),
    .Z(_04464_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _12459_ (.A1(_04463_),
    .A2(_04408_),
    .B(_04464_),
    .ZN(_04465_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _12460_ (.A1(_04319_),
    .A2(_04327_),
    .A3(_04380_),
    .ZN(_04466_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12461_ (.I(_04254_),
    .Z(_04467_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12462_ (.I(_04390_),
    .Z(_04468_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12463_ (.I(_04279_),
    .Z(_04469_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12464_ (.I(_04257_),
    .Z(_04470_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12465_ (.I(_04470_),
    .Z(_04471_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _12466_ (.A1(_04467_),
    .A2(_04468_),
    .B1(_04469_),
    .B2(_04471_),
    .ZN(_04472_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12467_ (.I(_04279_),
    .Z(_04473_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _12468_ (.A1(_04467_),
    .A2(_04471_),
    .A3(_04390_),
    .A4(_04473_),
    .ZN(_04474_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _12469_ (.A1(_04387_),
    .A2(_04472_),
    .B(_04474_),
    .ZN(_04475_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12470_ (.I(_04227_),
    .Z(_04476_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12471_ (.I(_04178_),
    .Z(_04477_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _12472_ (.A1(_04477_),
    .A2(_04476_),
    .ZN(_04478_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12473_ (.A1(_04236_),
    .A2(_04278_),
    .ZN(_04479_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12474_ (.I(_04385_),
    .Z(_04480_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12475_ (.A1(_04220_),
    .A2(_04480_),
    .ZN(_04481_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _12476_ (.A1(_04478_),
    .A2(_04479_),
    .A3(_04481_),
    .ZN(_04482_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12477_ (.I(_04404_),
    .Z(_04483_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _12478_ (.A1(_04174_),
    .A2(_04483_),
    .ZN(_04484_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12479_ (.I(_04267_),
    .Z(_04485_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12480_ (.A1(_04199_),
    .A2(_04485_),
    .ZN(_04486_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12481_ (.I(_04185_),
    .Z(_04487_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _12482_ (.A1(_03238_),
    .A2(_03182_),
    .A3(_04188_),
    .A4(_03410_),
    .ZN(_04488_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12483_ (.A1(_03413_),
    .A2(_04488_),
    .Z(_04489_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12484_ (.I(_04489_),
    .Z(_04490_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12485_ (.I(_04490_),
    .Z(_04491_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12486_ (.A1(_04487_),
    .A2(_04491_),
    .ZN(_04492_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _12487_ (.A1(_04484_),
    .A2(_04486_),
    .A3(_04492_),
    .ZN(_04493_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _12488_ (.A1(_04475_),
    .A2(_04482_),
    .A3(net71),
    .Z(_04494_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _12489_ (.A1(_04466_),
    .A2(_04494_),
    .Z(_04495_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _12490_ (.A1(_04462_),
    .A2(_04465_),
    .A3(_04495_),
    .ZN(_04496_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _12491_ (.A1(_04410_),
    .A2(_04412_),
    .Z(_04497_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12492_ (.I(_04416_),
    .Z(_04498_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _12493_ (.A1(_04292_),
    .A2(_04498_),
    .A3(_04423_),
    .ZN(_04499_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12494_ (.I(_04288_),
    .Z(_04500_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _12495_ (.A1(_04301_),
    .A2(_04500_),
    .A3(_04425_),
    .ZN(_04501_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12496_ (.A1(_04499_),
    .A2(_04501_),
    .Z(_04502_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12497_ (.A1(_04292_),
    .A2(_04288_),
    .ZN(_04503_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12498_ (.I(_04201_),
    .Z(_04504_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12499_ (.I(_04406_),
    .Z(_04505_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12500_ (.I(_04187_),
    .Z(_04506_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _12501_ (.A1(_04504_),
    .A2(_04206_),
    .B1(_04505_),
    .B2(_04506_),
    .ZN(_04507_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _12502_ (.A1(_04293_),
    .A2(_04504_),
    .A3(_04182_),
    .A4(_04505_),
    .ZN(_04508_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12503_ (.A1(_04398_),
    .A2(_04507_),
    .B(_04508_),
    .ZN(_04509_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12504_ (.I(_04396_),
    .Z(_04510_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12505_ (.I(_04510_),
    .Z(_04511_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12506_ (.I(_04511_),
    .Z(_04512_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12507_ (.A1(_04512_),
    .A2(_04302_),
    .ZN(_04513_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12508_ (.A1(_04509_),
    .A2(_04513_),
    .Z(_04514_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _12509_ (.A1(_04503_),
    .A2(_04514_),
    .Z(_04515_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _12510_ (.A1(_04497_),
    .A2(_04502_),
    .A3(_04515_),
    .Z(_04516_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _12511_ (.A1(_04440_),
    .A2(_04496_),
    .A3(_04516_),
    .Z(_04517_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _12512_ (.A1(_04438_),
    .A2(_04517_),
    .ZN(_04518_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _12513_ (.A1(_04435_),
    .A2(_04518_),
    .Z(_04519_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12514_ (.A1(_04431_),
    .A2(_04519_),
    .ZN(_04520_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _12515_ (.A1(_04223_),
    .A2(_04232_),
    .ZN(_04521_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12516_ (.I(net60),
    .Z(_04522_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _12517_ (.A1(_03333_),
    .A2(_04293_),
    .A3(_04522_),
    .ZN(_04523_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _12518_ (.A1(_03273_),
    .A2(_04243_),
    .A3(_04296_),
    .ZN(_04524_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12519_ (.I(_04266_),
    .Z(_04525_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _12520_ (.A1(_03317_),
    .A2(_04525_),
    .A3(_04164_),
    .Z(_04526_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _12521_ (.A1(_04523_),
    .A2(_04524_),
    .A3(_04526_),
    .ZN(_04527_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _12522_ (.A1(_04521_),
    .A2(_04527_),
    .ZN(_04528_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12523_ (.I(_04175_),
    .Z(_04529_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _12524_ (.A1(_03333_),
    .A2(_04529_),
    .A3(_04522_),
    .Z(_04530_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _12525_ (.A1(_04530_),
    .A2(_04193_),
    .A3(_04202_),
    .Z(_04531_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _12526_ (.A1(_04233_),
    .A2(_04245_),
    .A3(_04531_),
    .Z(_04532_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12527_ (.A1(_04532_),
    .A2(_04528_),
    .ZN(_04533_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _12528_ (.A1(_04172_),
    .A2(_04210_),
    .ZN(_04534_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12529_ (.I(_04333_),
    .Z(_04535_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12530_ (.A1(_04535_),
    .A2(_04171_),
    .ZN(_04536_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _12531_ (.A1(\filters.res_lut[1] ),
    .A2(_04168_),
    .ZN(_04537_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12532_ (.A1(_04523_),
    .A2(_04524_),
    .Z(_04538_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _12533_ (.A1(_04523_),
    .A2(_04524_),
    .Z(_04539_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _12534_ (.A1(_04537_),
    .A2(_04165_),
    .A3(_04538_),
    .B(_04539_),
    .ZN(_04540_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _12535_ (.A1(\filters.res_lut[2] ),
    .A2(_04169_),
    .ZN(_04541_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12536_ (.A1(_04165_),
    .A2(_04541_),
    .ZN(_04542_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12537_ (.A1(_04540_),
    .A2(_04542_),
    .Z(_04543_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12538_ (.A1(_04540_),
    .A2(_04542_),
    .Z(_04544_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _12539_ (.A1(_04536_),
    .A2(_04543_),
    .B(_04544_),
    .ZN(_04545_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _12540_ (.A1(_04172_),
    .A2(_04210_),
    .A3(_04533_),
    .Z(_04546_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _12541_ (.A1(_04545_),
    .A2(_04546_),
    .Z(_04547_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _12542_ (.A1(_04533_),
    .A2(_04534_),
    .B(_04547_),
    .ZN(_04548_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _12543_ (.A1(_04356_),
    .A2(_04249_),
    .A3(_04357_),
    .Z(_04549_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12544_ (.A1(_04545_),
    .A2(_04546_),
    .ZN(_04550_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _12545_ (.A1(_04549_),
    .A2(_04547_),
    .A3(_04550_),
    .ZN(_04551_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _12546_ (.A1(_04285_),
    .A2(_04213_),
    .A3(_04305_),
    .Z(_04552_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _12547_ (.A1(_04352_),
    .A2(_04359_),
    .A3(_04552_),
    .ZN(_04553_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12548_ (.A1(_04551_),
    .A2(_04553_),
    .ZN(_04554_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12549_ (.A1(_04551_),
    .A2(_04553_),
    .ZN(_04555_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _12550_ (.A1(_04548_),
    .A2(_04554_),
    .B(_04555_),
    .ZN(_04556_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _12551_ (.A1(_04362_),
    .A2(_04428_),
    .A3(_04309_),
    .Z(_04557_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _12552_ (.A1(_04556_),
    .A2(_04557_),
    .Z(_04558_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _12553_ (.A1(_04549_),
    .A2(_04545_),
    .A3(_04546_),
    .Z(_04559_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12554_ (.A1(_04528_),
    .A2(_04532_),
    .Z(_04560_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12555_ (.I(_04500_),
    .Z(_04561_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12556_ (.I(_04561_),
    .Z(_04562_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12557_ (.A1(_04468_),
    .A2(_04562_),
    .ZN(_04563_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12558_ (.A1(_04535_),
    .A2(_04537_),
    .ZN(_04564_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _12559_ (.A1(_03317_),
    .A2(_04506_),
    .A3(_04164_),
    .ZN(_04565_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12560_ (.I(_04226_),
    .Z(_04566_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _12561_ (.A1(_03255_),
    .A2(_04566_),
    .A3(_04504_),
    .ZN(_04567_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12562_ (.A1(_04565_),
    .A2(_04567_),
    .ZN(_04568_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12563_ (.A1(_04565_),
    .A2(_04567_),
    .ZN(_04569_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _12564_ (.A1(_04564_),
    .A2(_04568_),
    .B(_04569_),
    .ZN(_04570_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12565_ (.A1(_04297_),
    .A2(_04498_),
    .ZN(_04571_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _12566_ (.A1(_04570_),
    .A2(_04571_),
    .ZN(_04572_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _12567_ (.A1(_04570_),
    .A2(_04571_),
    .Z(_04573_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _12568_ (.A1(_04563_),
    .A2(_04572_),
    .B(_04573_),
    .ZN(_04574_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12569_ (.I(_04231_),
    .Z(_04575_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12570_ (.I(_04575_),
    .Z(_04576_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12571_ (.A1(_04354_),
    .A2(_04576_),
    .ZN(_04577_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12572_ (.I(_04525_),
    .Z(_04578_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _12573_ (.A1(_03302_),
    .A2(_04332_),
    .A3(_04578_),
    .ZN(_04579_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _12574_ (.A1(_04565_),
    .A2(_04567_),
    .A3(_04579_),
    .Z(_04580_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12575_ (.A1(_04577_),
    .A2(_04580_),
    .ZN(_04581_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12576_ (.A1(_04521_),
    .A2(_04527_),
    .Z(_04582_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12577_ (.A1(_04581_),
    .A2(_04582_),
    .Z(_04583_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _12578_ (.A1(_04540_),
    .A2(_04542_),
    .A3(_04536_),
    .Z(_04584_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12579_ (.A1(_04583_),
    .A2(_04584_),
    .Z(_04585_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _12580_ (.A1(_04574_),
    .A2(_04585_),
    .Z(_04586_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _12581_ (.A1(_04559_),
    .A2(_04560_),
    .A3(_04586_),
    .Z(_04587_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12582_ (.A1(_04574_),
    .A2(_04585_),
    .Z(_04588_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _12583_ (.A1(_04583_),
    .A2(_04584_),
    .B(_04588_),
    .ZN(_04589_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _12584_ (.A1(_04560_),
    .A2(_04586_),
    .B(_04559_),
    .ZN(_04590_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _12585_ (.A1(_04587_),
    .A2(_04589_),
    .A3(_04590_),
    .Z(_04591_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12586_ (.A1(_04581_),
    .A2(_04582_),
    .Z(_04592_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12587_ (.A1(_03272_),
    .A2(_04242_),
    .ZN(_04593_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12588_ (.I(_04593_),
    .Z(_04594_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12589_ (.A1(_04594_),
    .A2(_04171_),
    .ZN(_04595_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12590_ (.I(_04529_),
    .Z(_04596_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12591_ (.I(_04596_),
    .Z(_04597_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12592_ (.A1(_04468_),
    .A2(_04597_),
    .ZN(_04598_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12593_ (.I(_04506_),
    .Z(_04599_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12594_ (.I(_04296_),
    .Z(_04600_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12595_ (.I(_04600_),
    .Z(_04601_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _12596_ (.A1(_04297_),
    .A2(_04599_),
    .B1(_04601_),
    .B2(_04353_),
    .ZN(_04602_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _12597_ (.A1(_04353_),
    .A2(_04297_),
    .A3(_04599_),
    .A4(_04601_),
    .ZN(_04603_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12598_ (.A1(_04598_),
    .A2(_04602_),
    .B(_04603_),
    .ZN(_04604_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12599_ (.A1(_04261_),
    .A2(_04541_),
    .ZN(_04605_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _12600_ (.A1(_04604_),
    .A2(_04605_),
    .Z(_04606_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12601_ (.A1(_04604_),
    .A2(_04605_),
    .Z(_04607_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _12602_ (.A1(_04595_),
    .A2(_04606_),
    .B(_04607_),
    .ZN(_04608_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _12603_ (.A1(_04563_),
    .A2(_04572_),
    .ZN(_04609_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _12604_ (.A1(_04592_),
    .A2(_04608_),
    .A3(_04609_),
    .Z(_04610_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12605_ (.A1(_04577_),
    .A2(_04580_),
    .Z(_04611_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _12606_ (.I(_04611_),
    .ZN(_04612_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _12607_ (.A1(_03256_),
    .A2(_04566_),
    .ZN(_04613_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12608_ (.A1(_04613_),
    .A2(_04171_),
    .ZN(_04614_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12609_ (.I(_04369_),
    .Z(_04615_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12610_ (.I(_04578_),
    .Z(_04616_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12611_ (.I(_04599_),
    .Z(_04617_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _12612_ (.A1(_04615_),
    .A2(_04468_),
    .A3(_04616_),
    .A4(_04617_),
    .ZN(_04618_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12613_ (.I(_04498_),
    .Z(_04619_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12614_ (.A1(_04615_),
    .A2(_04619_),
    .ZN(_04620_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12615_ (.A1(_04618_),
    .A2(_04620_),
    .ZN(_04621_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12616_ (.A1(_04541_),
    .A2(_04618_),
    .ZN(_04622_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _12617_ (.A1(_04614_),
    .A2(_04621_),
    .B(_04622_),
    .ZN(_04623_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _12618_ (.A1(_04604_),
    .A2(_04605_),
    .A3(_04595_),
    .ZN(_04624_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12619_ (.A1(_04623_),
    .A2(_04624_),
    .Z(_04625_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _12620_ (.A1(_04623_),
    .A2(_04624_),
    .Z(_04626_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _12621_ (.A1(_04612_),
    .A2(_04625_),
    .B(_04626_),
    .ZN(_04627_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12622_ (.I(_04354_),
    .Z(_04628_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12623_ (.I(_04420_),
    .Z(_04629_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12624_ (.I(_04629_),
    .Z(_04630_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12625_ (.I(_04630_),
    .Z(_04631_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _12626_ (.I(_04619_),
    .Z(_04632_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12627_ (.I(_04616_),
    .Z(_04633_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12628_ (.I(_04617_),
    .Z(_04634_));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 _12629_ (.A1(_03256_),
    .A2(_04566_),
    .A3(_04633_),
    .A4(_04634_),
    .Z(_04635_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _12630_ (.A1(_04615_),
    .A2(_04632_),
    .A3(_04635_),
    .ZN(_04636_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _12631_ (.A1(_03256_),
    .A2(_04566_),
    .A3(_04633_),
    .A4(_04634_),
    .ZN(_04637_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_4 _12632_ (.A1(_04613_),
    .A2(_04541_),
    .B1(_04637_),
    .B2(_04594_),
    .ZN(_04638_));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 _12633_ (.A1(_04628_),
    .A2(_04631_),
    .A3(_04636_),
    .A4(_04638_),
    .Z(_04639_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _12634_ (.A1(_04628_),
    .A2(_04631_),
    .B1(_04636_),
    .B2(_04638_),
    .ZN(_04640_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12635_ (.I(_04207_),
    .Z(_04641_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12636_ (.I(_04641_),
    .Z(_04642_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12637_ (.I(_04642_),
    .Z(_04643_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _12638_ (.I(_04643_),
    .Z(_04644_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12639_ (.I(_04644_),
    .Z(_04645_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _12640_ (.A1(_04628_),
    .A2(_04645_),
    .A3(_04635_),
    .ZN(_04646_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _12641_ (.A1(_04639_),
    .A2(_04640_),
    .B(_04646_),
    .ZN(_04647_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12642_ (.A1(\filters.res_lut[0] ),
    .A2(_04170_),
    .ZN(_04648_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _12643_ (.A1(_04594_),
    .A2(_04537_),
    .B1(_04648_),
    .B2(_04261_),
    .ZN(_04649_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12644_ (.A1(_04618_),
    .A2(_04649_),
    .ZN(_04650_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _12645_ (.A1(_04639_),
    .A2(_04640_),
    .A3(_04646_),
    .B(_04650_),
    .ZN(_04651_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12646_ (.A1(_04647_),
    .A2(_04651_),
    .ZN(_04652_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12647_ (.A1(_04535_),
    .A2(_04648_),
    .ZN(_04653_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12648_ (.A1(_04354_),
    .A2(_04601_),
    .ZN(_04654_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _12649_ (.A1(_04653_),
    .A2(_04654_),
    .A3(_04598_),
    .Z(_04655_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12650_ (.I0(_04644_),
    .I1(_04620_),
    .S(_04618_),
    .Z(_04656_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _12651_ (.A1(_04614_),
    .A2(_04656_),
    .ZN(_04657_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _12652_ (.I(_04636_),
    .ZN(_04658_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _12653_ (.A1(_04658_),
    .A2(_04639_),
    .Z(_04659_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _12654_ (.A1(_04655_),
    .A2(_04657_),
    .A3(_04659_),
    .ZN(_04660_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _12655_ (.A1(_04623_),
    .A2(_04624_),
    .A3(_04612_),
    .Z(_04661_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _12656_ (.A1(_04652_),
    .A2(_04660_),
    .B(_04661_),
    .ZN(_04662_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _12657_ (.A1(_04655_),
    .A2(_04657_),
    .A3(_04659_),
    .ZN(_04663_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _12658_ (.A1(_04639_),
    .A2(_04640_),
    .B(_04646_),
    .C(_04650_),
    .ZN(_04664_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _12659_ (.A1(_04322_),
    .A2(_04633_),
    .B1(_04634_),
    .B2(_04615_),
    .ZN(_04665_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12660_ (.A1(_04594_),
    .A2(_04637_),
    .B(_04628_),
    .ZN(_04666_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12661_ (.I(_04632_),
    .Z(_04667_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12662_ (.A1(_04667_),
    .A2(_04635_),
    .B(_04646_),
    .ZN(_04668_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _12663_ (.A1(_04665_),
    .A2(_04666_),
    .A3(_04668_),
    .ZN(_04669_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _12664_ (.A1(_04647_),
    .A2(_04651_),
    .B1(_04664_),
    .B2(_04669_),
    .ZN(_04670_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _12665_ (.A1(_04657_),
    .A2(_04659_),
    .B(_04655_),
    .ZN(_04671_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12666_ (.A1(_04657_),
    .A2(_04659_),
    .ZN(_04672_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _12667_ (.A1(_04663_),
    .A2(_04670_),
    .B(_04671_),
    .C(_04672_),
    .ZN(_04673_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _12668_ (.A1(_04610_),
    .A2(_04627_),
    .B1(_04662_),
    .B2(_04673_),
    .ZN(_04674_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _12669_ (.A1(_04610_),
    .A2(_04627_),
    .ZN(_04675_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _12670_ (.I(_04560_),
    .ZN(_04676_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12671_ (.A1(_04676_),
    .A2(_04586_),
    .Z(_04677_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _12672_ (.A1(_04674_),
    .A2(_04675_),
    .B(_04677_),
    .ZN(_04678_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12673_ (.A1(_04608_),
    .A2(_04609_),
    .ZN(_04679_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12674_ (.A1(_04608_),
    .A2(_04609_),
    .ZN(_04680_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _12675_ (.A1(_04592_),
    .A2(_04679_),
    .B(_04680_),
    .ZN(_04681_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _12676_ (.A1(_04677_),
    .A2(_04674_),
    .A3(_04675_),
    .B(_04681_),
    .ZN(_04682_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _12677_ (.A1(_04587_),
    .A2(_04590_),
    .B(_04589_),
    .ZN(_04683_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _12678_ (.A1(_04591_),
    .A2(_04678_),
    .A3(_04682_),
    .A4(_04683_),
    .ZN(_04684_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _12679_ (.A1(_04551_),
    .A2(_04553_),
    .A3(_04548_),
    .Z(_04685_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _12680_ (.A1(_04559_),
    .A2(_04560_),
    .A3(_04586_),
    .ZN(_04686_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12681_ (.A1(_04589_),
    .A2(_04590_),
    .B(_04686_),
    .ZN(_04687_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _12682_ (.A1(_04687_),
    .A2(_04685_),
    .ZN(_04688_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _12683_ (.A1(_04685_),
    .A2(_04687_),
    .ZN(_04689_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _12684_ (.A1(_04684_),
    .A2(_04688_),
    .B(_04689_),
    .ZN(_04690_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _12685_ (.A1(_04556_),
    .A2(_04557_),
    .ZN(_04691_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _12686_ (.A1(_04431_),
    .A2(_04519_),
    .B1(_04558_),
    .B2(_04690_),
    .C(_04691_),
    .ZN(_04692_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _12687_ (.A1(_04520_),
    .A2(_04692_),
    .Z(_04693_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12688_ (.I(_04467_),
    .Z(_04694_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12689_ (.I(_04385_),
    .Z(_04695_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12690_ (.I(_04695_),
    .Z(_04696_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12691_ (.I(_04392_),
    .Z(_04697_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _12692_ (.A1(_04694_),
    .A2(_04281_),
    .B1(_04696_),
    .B2(_04697_),
    .ZN(_04698_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12693_ (.I(_04255_),
    .Z(_04699_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _12694_ (.A1(_04699_),
    .A2(_04697_),
    .A3(_04469_),
    .A4(_04696_),
    .ZN(_04700_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _12695_ (.A1(_04478_),
    .A2(_04698_),
    .B(_04700_),
    .ZN(_04701_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12696_ (.A1(_04388_),
    .A2(_04480_),
    .ZN(_04702_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12697_ (.I(_04257_),
    .Z(_04703_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12698_ (.A1(_04703_),
    .A2(_04180_),
    .ZN(_04704_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12699_ (.I(_04476_),
    .Z(_04705_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12700_ (.A1(_04705_),
    .A2(_04268_),
    .ZN(_04706_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _12701_ (.A1(_04702_),
    .A2(_04704_),
    .A3(_04706_),
    .ZN(_04707_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12702_ (.A1(_04701_),
    .A2(_04707_),
    .ZN(_04708_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12703_ (.A1(_04265_),
    .A2(_04491_),
    .ZN(_04709_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12704_ (.I(_03184_),
    .Z(_04710_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12705_ (.I0(\filters.high[12] ),
    .I1(\filters.band[12] ),
    .S(_04710_),
    .Z(_04711_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12706_ (.I(_04711_),
    .Z(_04712_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12707_ (.I(_04712_),
    .Z(_04713_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _12708_ (.A1(_04186_),
    .A2(_04713_),
    .ZN(_04714_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12709_ (.A1(_04274_),
    .A2(_04295_),
    .ZN(_04715_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _12710_ (.A1(_04709_),
    .A2(_04714_),
    .A3(_04715_),
    .ZN(_04716_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _12711_ (.I(_04716_),
    .ZN(_04717_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12712_ (.A1(_04701_),
    .A2(_04707_),
    .ZN(_04718_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12713_ (.A1(_04708_),
    .A2(_04717_),
    .B(_04718_),
    .ZN(_04719_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12714_ (.A1(_04366_),
    .A2(_04279_),
    .Z(_04720_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _12715_ (.A1(_03271_),
    .A2(_04241_),
    .A3(_04376_),
    .Z(_04721_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _12716_ (.A1(_03288_),
    .A2(_04316_),
    .A3(_04197_),
    .Z(_04722_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _12717_ (.A1(_04720_),
    .A2(_04721_),
    .A3(_04722_),
    .ZN(_04723_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12718_ (.A1(_04458_),
    .A2(_04459_),
    .ZN(_04724_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12719_ (.A1(_04458_),
    .A2(_04459_),
    .ZN(_04725_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _12720_ (.A1(_04457_),
    .A2(_04724_),
    .B(_04725_),
    .ZN(_04726_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12721_ (.A1(_04723_),
    .A2(_04726_),
    .ZN(_04727_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12722_ (.I(_04236_),
    .Z(_04728_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _12723_ (.I(_04477_),
    .Z(_04729_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _12724_ (.A1(_04728_),
    .A2(_04695_),
    .B1(_04729_),
    .B2(_04259_),
    .ZN(_04730_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _12725_ (.A1(_04728_),
    .A2(_04259_),
    .A3(_04695_),
    .A4(_04729_),
    .ZN(_04731_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _12726_ (.A1(_04706_),
    .A2(_04730_),
    .B(_04731_),
    .ZN(_04732_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12727_ (.A1(_04228_),
    .A2(_04272_),
    .ZN(_04733_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12728_ (.A1(_04253_),
    .A2(_04179_),
    .ZN(_04734_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12729_ (.A1(_04258_),
    .A2(_04485_),
    .ZN(_04735_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _12730_ (.A1(_04733_),
    .A2(_04734_),
    .A3(_04735_),
    .ZN(_04736_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12731_ (.I(_04711_),
    .Z(_04737_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12732_ (.A1(_04173_),
    .A2(_04737_),
    .ZN(_04738_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12733_ (.I0(\filters.high[13] ),
    .I1(\filters.band[13] ),
    .S(_04710_),
    .Z(_04739_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12734_ (.I(_04739_),
    .Z(_04740_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12735_ (.A1(_04184_),
    .A2(_04740_),
    .ZN(_04741_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12736_ (.I(_04198_),
    .Z(_04742_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12737_ (.A1(_04510_),
    .A2(_04742_),
    .ZN(_04743_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _12738_ (.A1(_04738_),
    .A2(_04741_),
    .A3(_04743_),
    .ZN(_04744_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _12739_ (.A1(_04732_),
    .A2(_04736_),
    .A3(_04744_),
    .Z(_04745_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12740_ (.A1(_04727_),
    .A2(_04745_),
    .Z(_04746_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12741_ (.A1(_04727_),
    .A2(_04745_),
    .Z(_04747_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _12742_ (.A1(_04719_),
    .A2(_04746_),
    .B(_04747_),
    .ZN(_04748_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _12743_ (.I(_04748_),
    .ZN(_04749_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12744_ (.I(_04489_),
    .Z(_04750_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12745_ (.I(_04750_),
    .Z(_04751_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12746_ (.I(_04751_),
    .Z(_04752_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12747_ (.I(_04752_),
    .Z(_04753_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12748_ (.A1(_04286_),
    .A2(_04753_),
    .ZN(_04754_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12749_ (.A1(_04741_),
    .A2(_04743_),
    .Z(_04755_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _12750_ (.A1(_04741_),
    .A2(_04743_),
    .Z(_04756_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12751_ (.A1(_04738_),
    .A2(_04755_),
    .B(_04756_),
    .ZN(_04757_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12752_ (.I(_04713_),
    .Z(_04758_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12753_ (.I(_04758_),
    .Z(_04759_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12754_ (.A1(_04641_),
    .A2(_04759_),
    .ZN(_04760_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _12755_ (.A1(_04754_),
    .A2(_04757_),
    .A3(_04760_),
    .Z(_04761_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12756_ (.A1(_04749_),
    .A2(_04761_),
    .ZN(_04762_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12757_ (.A1(_04287_),
    .A2(_04505_),
    .ZN(_04763_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12758_ (.I(_04211_),
    .Z(_04764_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12759_ (.I(_04764_),
    .Z(_04765_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12760_ (.I(_04753_),
    .Z(_04766_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12761_ (.A1(_04714_),
    .A2(_04715_),
    .Z(_04767_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _12762_ (.A1(_04714_),
    .A2(_04715_),
    .Z(_04768_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12763_ (.A1(_04709_),
    .A2(_04767_),
    .B(_04768_),
    .ZN(_04769_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _12764_ (.A1(_04765_),
    .A2(_04766_),
    .B(_04769_),
    .ZN(_04770_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _12765_ (.A1(_04765_),
    .A2(_04766_),
    .A3(_04769_),
    .ZN(_04771_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12766_ (.A1(_04763_),
    .A2(_04770_),
    .B(_04771_),
    .ZN(_04772_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _12767_ (.A1(_04748_),
    .A2(_04761_),
    .ZN(_04773_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12768_ (.A1(_04772_),
    .A2(_04773_),
    .ZN(_04774_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12769_ (.A1(_04762_),
    .A2(_04774_),
    .ZN(_04775_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12770_ (.I(_04442_),
    .Z(_04776_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12771_ (.A1(\filters.cutoff_lut[11] ),
    .A2(_04776_),
    .ZN(_04777_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _12772_ (.A1(_04593_),
    .A2(_04777_),
    .ZN(_04778_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12773_ (.A1(\filters.cutoff_lut[13] ),
    .A2(_04442_),
    .Z(_04779_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12774_ (.I(_04779_),
    .Z(_04780_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12775_ (.I(_04780_),
    .Z(_04781_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _12776_ (.A1(_03200_),
    .A2(_04216_),
    .A3(_04781_),
    .ZN(_04782_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12777_ (.A1(\filters.cutoff_lut[12] ),
    .A2(_04442_),
    .Z(_04783_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12778_ (.I(_04783_),
    .Z(_04784_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _12779_ (.A1(_03253_),
    .A2(_04225_),
    .A3(_04784_),
    .ZN(_04785_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _12780_ (.A1(_04782_),
    .A2(_04785_),
    .Z(_04786_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _12781_ (.A1(_04778_),
    .A2(_04786_),
    .ZN(_04787_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _12782_ (.A1(_04721_),
    .A2(_04722_),
    .Z(_04788_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12783_ (.A1(_04721_),
    .A2(_04722_),
    .Z(_04789_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _12784_ (.A1(_04720_),
    .A2(_04788_),
    .B(_04789_),
    .ZN(_04790_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12785_ (.I(_04783_),
    .Z(_04791_));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 _12786_ (.A1(_04311_),
    .A2(_04321_),
    .A3(_04444_),
    .A4(_04791_),
    .Z(_04792_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _12787_ (.A1(_03315_),
    .A2(_04323_),
    .A3(net59),
    .ZN(_04793_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _12788_ (.A1(net63),
    .A2(_04195_),
    .A3(_04374_),
    .ZN(_04794_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _12789_ (.A1(_03301_),
    .A2(_04314_),
    .A3(_04276_),
    .ZN(_04795_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _12790_ (.A1(_04793_),
    .A2(_04794_),
    .A3(_04795_),
    .ZN(_04796_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _12791_ (.A1(_04792_),
    .A2(_04796_),
    .ZN(_04797_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _12792_ (.A1(_04790_),
    .A2(_04797_),
    .ZN(_04798_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12793_ (.A1(_04787_),
    .A2(_04798_),
    .Z(_04799_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12794_ (.I(_04443_),
    .Z(_04800_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12795_ (.I(_04800_),
    .Z(_04801_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12796_ (.I(_04801_),
    .Z(_04802_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12797_ (.I(_04783_),
    .Z(_04803_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12798_ (.I(_04803_),
    .Z(_04804_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12799_ (.I(_04804_),
    .Z(_04805_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12800_ (.I(_04805_),
    .Z(_04806_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _12801_ (.A1(_04322_),
    .A2(_04802_),
    .B1(_04806_),
    .B2(_04313_),
    .ZN(_04807_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _12802_ (.A1(_04792_),
    .A2(_04807_),
    .ZN(_04808_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _12803_ (.A1(_04723_),
    .A2(_04726_),
    .Z(_04809_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12804_ (.A1(_04808_),
    .A2(_04809_),
    .ZN(_04810_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12805_ (.A1(_04799_),
    .A2(_04810_),
    .Z(_04811_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _12806_ (.A1(_04746_),
    .A2(_04719_),
    .ZN(_04812_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _12807_ (.A1(_04799_),
    .A2(_04808_),
    .A3(_04809_),
    .ZN(_04813_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _12808_ (.A1(_04811_),
    .A2(net50),
    .B(_04813_),
    .ZN(_04814_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12809_ (.A1(_04787_),
    .A2(_04798_),
    .ZN(_04815_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _12810_ (.A1(\filters.cutoff_lut[14] ),
    .A2(_04441_),
    .Z(_04816_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12811_ (.I(_04816_),
    .Z(_04817_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12812_ (.I(_04817_),
    .Z(_04818_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12813_ (.I(_04818_),
    .Z(_04819_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12814_ (.I(_04819_),
    .Z(_04820_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _12815_ (.A1(_04313_),
    .A2(_04820_),
    .ZN(_04821_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _12816_ (.A1(_03287_),
    .A2(_04197_),
    .A3(_04444_),
    .ZN(_04822_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _12817_ (.A1(_03271_),
    .A2(_04242_),
    .A3(_04784_),
    .ZN(_04823_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12818_ (.I(_04780_),
    .Z(_04824_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12819_ (.I(_04824_),
    .Z(_04825_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _12820_ (.A1(_03254_),
    .A2(_04225_),
    .A3(_04825_),
    .ZN(_04826_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _12821_ (.A1(_04822_),
    .A2(_04823_),
    .A3(_04826_),
    .Z(_04827_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _12822_ (.A1(_04821_),
    .A2(_04827_),
    .ZN(_04828_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12823_ (.A1(_04794_),
    .A2(_04795_),
    .Z(_04829_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _12824_ (.A1(_04794_),
    .A2(_04795_),
    .Z(_04830_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _12825_ (.A1(_04793_),
    .A2(_04829_),
    .B(_04830_),
    .ZN(_04831_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12826_ (.A1(_04782_),
    .A2(_04785_),
    .ZN(_04832_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _12827_ (.A1(_04778_),
    .A2(_04786_),
    .B(_04832_),
    .ZN(_04833_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _12828_ (.A1(_04324_),
    .A2(_04729_),
    .ZN(_04834_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12829_ (.A1(_04316_),
    .A2(_04480_),
    .ZN(_04835_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12830_ (.A1(_04473_),
    .A2(_04377_),
    .ZN(_04836_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _12831_ (.A1(_04834_),
    .A2(_04835_),
    .A3(_04836_),
    .Z(_04837_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _12832_ (.A1(_04831_),
    .A2(_04833_),
    .A3(_04837_),
    .ZN(_04838_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12833_ (.A1(_04828_),
    .A2(_04838_),
    .Z(_04839_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12834_ (.A1(_04815_),
    .A2(_04839_),
    .Z(_04840_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12835_ (.A1(_04732_),
    .A2(_04736_),
    .ZN(_04841_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _12836_ (.I(_04744_),
    .ZN(_04842_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12837_ (.A1(_04732_),
    .A2(_04736_),
    .ZN(_04843_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _12838_ (.A1(_04841_),
    .A2(_04842_),
    .B(_04843_),
    .ZN(_04844_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12839_ (.A1(_04792_),
    .A2(_04796_),
    .ZN(_04845_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _12840_ (.A1(_04790_),
    .A2(_04797_),
    .B(_04845_),
    .ZN(_04846_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12841_ (.I(_04220_),
    .Z(_04847_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _12842_ (.I(_04237_),
    .Z(_04848_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _12843_ (.A1(_04847_),
    .A2(_04269_),
    .B1(_04181_),
    .B2(_04848_),
    .ZN(_04849_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12844_ (.I(_04703_),
    .Z(_04850_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _12845_ (.A1(_04848_),
    .A2(_04850_),
    .A3(_04268_),
    .A4(_04181_),
    .ZN(_04851_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _12846_ (.A1(_04733_),
    .A2(_04849_),
    .B(_04851_),
    .ZN(_04852_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _12847_ (.A1(_04476_),
    .A2(_04396_),
    .Z(_04853_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12848_ (.I(_04271_),
    .Z(_04854_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _12849_ (.A1(_03364_),
    .A2(_04219_),
    .A3(_04854_),
    .ZN(_04855_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _12850_ (.A1(_03349_),
    .A2(net68),
    .A3(_04192_),
    .ZN(_04856_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _12851_ (.A1(_04853_),
    .A2(_04855_),
    .A3(_04856_),
    .Z(_04857_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12852_ (.I(_04739_),
    .Z(_04858_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12853_ (.A1(_04174_),
    .A2(_04858_),
    .ZN(_04859_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12854_ (.I0(\filters.high[14] ),
    .I1(\filters.band[14] ),
    .S(_04710_),
    .Z(_04860_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12855_ (.I(_04860_),
    .Z(_04861_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12856_ (.I(_04861_),
    .Z(_04862_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _12857_ (.A1(_04400_),
    .A2(_04862_),
    .ZN(_04863_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12858_ (.I(_04483_),
    .Z(_04864_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12859_ (.A1(_04200_),
    .A2(_04864_),
    .ZN(_04865_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _12860_ (.A1(_04859_),
    .A2(_04863_),
    .A3(_04865_),
    .ZN(_04866_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _12861_ (.A1(_04852_),
    .A2(_04857_),
    .A3(_04866_),
    .Z(_04867_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12862_ (.A1(_04867_),
    .A2(_04846_),
    .Z(_04868_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12863_ (.A1(_04868_),
    .A2(_04844_),
    .Z(_04869_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _12864_ (.A1(_04840_),
    .A2(_04869_),
    .Z(_04870_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12865_ (.A1(_04814_),
    .A2(_04870_),
    .ZN(_04871_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _12866_ (.A1(_04772_),
    .A2(_04773_),
    .ZN(_04872_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12867_ (.A1(_04814_),
    .A2(_04870_),
    .ZN(_04873_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12868_ (.A1(_04871_),
    .A2(_04872_),
    .B(_04873_),
    .ZN(_04874_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12869_ (.A1(_04815_),
    .A2(_04839_),
    .Z(_04875_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _12870_ (.A1(_04840_),
    .A2(_04869_),
    .B(_04875_),
    .ZN(_04876_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _12871_ (.A1(_04828_),
    .A2(_04838_),
    .ZN(_04877_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _12872_ (.A1(_04821_),
    .A2(_04827_),
    .ZN(_04878_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _12873_ (.A1(\filters.cutoff_lut[15] ),
    .A2(_04441_),
    .Z(_04879_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12874_ (.I(_04879_),
    .Z(_04880_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _12875_ (.I(_04880_),
    .Z(_04881_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12876_ (.I(_04881_),
    .Z(_04882_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _12877_ (.A1(_03199_),
    .A2(_04215_),
    .A3(_04882_),
    .ZN(_04883_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12878_ (.I(_04816_),
    .Z(_04884_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _12879_ (.A1(_03253_),
    .A2(_04224_),
    .A3(_04884_),
    .ZN(_04885_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _12880_ (.A1(_04883_),
    .A2(_04885_),
    .ZN(_04886_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _12881_ (.A1(_03302_),
    .A2(_04332_),
    .A3(_04800_),
    .ZN(_04887_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _12882_ (.A1(_03287_),
    .A2(_04196_),
    .A3(_04803_),
    .ZN(_04888_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _12883_ (.A1(_03272_),
    .A2(_04242_),
    .A3(_04824_),
    .ZN(_04889_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _12884_ (.A1(_04887_),
    .A2(_04888_),
    .A3(_04889_),
    .Z(_04890_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12885_ (.A1(_04886_),
    .A2(_04890_),
    .Z(_04891_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _12886_ (.A1(_04449_),
    .A2(_04696_),
    .B1(_04378_),
    .B2(_04469_),
    .ZN(_04892_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12887_ (.I(_04316_),
    .Z(_04893_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _12888_ (.A1(_04893_),
    .A2(_04469_),
    .A3(_04696_),
    .A4(_04378_),
    .ZN(_04894_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _12889_ (.A1(_04834_),
    .A2(_04892_),
    .B(_04894_),
    .ZN(_04895_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12890_ (.I(_04777_),
    .Z(_04896_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _12891_ (.A1(_04261_),
    .A2(_04896_),
    .ZN(_04897_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12892_ (.A1(_04823_),
    .A2(_04826_),
    .ZN(_04898_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12893_ (.A1(_04823_),
    .A2(_04826_),
    .ZN(_04899_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _12894_ (.A1(_04897_),
    .A2(_04898_),
    .B(_04899_),
    .ZN(_04900_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12895_ (.A1(_04367_),
    .A2(_04268_),
    .ZN(_04901_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _12896_ (.A1(_03332_),
    .A2(_04371_),
    .A3(net60),
    .ZN(_04902_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _12897_ (.A1(_03316_),
    .A2(_04163_),
    .A3(_04450_),
    .ZN(_04903_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _12898_ (.A1(_04902_),
    .A2(_04903_),
    .ZN(_04904_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _12899_ (.A1(_04901_),
    .A2(_04904_),
    .ZN(_04905_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _12900_ (.A1(_04895_),
    .A2(_04900_),
    .A3(_04905_),
    .ZN(_04906_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _12901_ (.A1(_04878_),
    .A2(_04891_),
    .A3(_04906_),
    .ZN(_04907_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12902_ (.A1(_04852_),
    .A2(_04857_),
    .ZN(_04908_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _12903_ (.I(_04866_),
    .ZN(_04909_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12904_ (.A1(_04852_),
    .A2(_04857_),
    .ZN(_04910_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12905_ (.A1(_04908_),
    .A2(_04909_),
    .B(_04910_),
    .ZN(_04911_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12906_ (.A1(_04833_),
    .A2(_04837_),
    .ZN(_04912_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12907_ (.A1(_04833_),
    .A2(_04837_),
    .ZN(_04913_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _12908_ (.A1(_04831_),
    .A2(_04912_),
    .B(_04913_),
    .ZN(_04914_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12909_ (.A1(_04855_),
    .A2(_04856_),
    .ZN(_04915_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12910_ (.A1(_04855_),
    .A2(_04856_),
    .ZN(_04916_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _12911_ (.A1(_04853_),
    .A2(_04915_),
    .B(_04916_),
    .ZN(_04917_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _12912_ (.A1(_04229_),
    .A2(_04483_),
    .ZN(_04918_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12913_ (.A1(_04470_),
    .A2(_04510_),
    .ZN(_04919_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12914_ (.A1(_04237_),
    .A2(_04273_),
    .ZN(_04920_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _12915_ (.A1(_04918_),
    .A2(_04919_),
    .A3(_04920_),
    .Z(_04921_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _12916_ (.A1(_04921_),
    .A2(_04917_),
    .ZN(_04922_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12917_ (.I(_04861_),
    .Z(_04923_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12918_ (.I(_04923_),
    .Z(_04924_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12919_ (.A1(_04175_),
    .A2(_04924_),
    .ZN(_04925_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12920_ (.I0(\filters.high[15] ),
    .I1(\filters.band[15] ),
    .S(_03185_),
    .Z(_04926_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12921_ (.I(_04926_),
    .Z(_04927_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12922_ (.A1(_04487_),
    .A2(_04927_),
    .ZN(_04928_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12923_ (.I(_04491_),
    .Z(_04929_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12924_ (.A1(_04295_),
    .A2(_04929_),
    .ZN(_04930_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _12925_ (.A1(_04925_),
    .A2(_04928_),
    .A3(_04930_),
    .Z(_04931_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _12926_ (.A1(_04922_),
    .A2(_04931_),
    .ZN(_04932_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _12927_ (.A1(_04911_),
    .A2(_04914_),
    .A3(_04932_),
    .ZN(_04933_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _12928_ (.A1(_04877_),
    .A2(_04907_),
    .A3(_04933_),
    .Z(_04934_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _12929_ (.A1(_04876_),
    .A2(_04934_),
    .ZN(_04935_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _12930_ (.A1(_04632_),
    .A2(_04759_),
    .B(_04757_),
    .ZN(_04936_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _12931_ (.A1(_04644_),
    .A2(_04759_),
    .A3(_04757_),
    .ZN(_04937_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _12932_ (.A1(_04754_),
    .A2(_04936_),
    .B(_04937_),
    .ZN(_04938_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12933_ (.A1(_04846_),
    .A2(_04867_),
    .Z(_04939_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _12934_ (.A1(_04844_),
    .A2(_04868_),
    .B(_04939_),
    .ZN(_04940_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12935_ (.A1(_04287_),
    .A2(_04759_),
    .ZN(_04941_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12936_ (.A1(_04863_),
    .A2(_04865_),
    .Z(_04942_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _12937_ (.A1(_04863_),
    .A2(_04865_),
    .Z(_04943_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _12938_ (.A1(_04859_),
    .A2(_04942_),
    .B(_04943_),
    .ZN(_04944_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12939_ (.I(_04858_),
    .Z(_04945_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12940_ (.I(_04945_),
    .Z(_04946_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12941_ (.A1(_04416_),
    .A2(_04946_),
    .ZN(_04947_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _12942_ (.A1(_04941_),
    .A2(_04944_),
    .A3(_04947_),
    .Z(_04948_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _12943_ (.A1(_04940_),
    .A2(_04948_),
    .ZN(_04949_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _12944_ (.A1(_04938_),
    .A2(_04949_),
    .ZN(_04950_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12945_ (.A1(_04935_),
    .A2(_04950_),
    .Z(_04951_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _12946_ (.A1(_04775_),
    .A2(_04874_),
    .A3(_04951_),
    .ZN(_04952_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12947_ (.A1(_04475_),
    .A2(_04482_),
    .ZN(_04953_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _12948_ (.I(_04493_),
    .ZN(_04954_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12949_ (.A1(_04475_),
    .A2(_04482_),
    .ZN(_04955_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _12950_ (.A1(_04953_),
    .A2(_04954_),
    .B(_04955_),
    .ZN(_04956_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12951_ (.A1(_04456_),
    .A2(_04460_),
    .Z(_04957_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _12952_ (.A1(_04701_),
    .A2(_04707_),
    .A3(_04716_),
    .Z(_04958_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _12953_ (.A1(_04957_),
    .A2(_04958_),
    .Z(_04959_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12954_ (.A1(_04957_),
    .A2(_04958_),
    .Z(_04960_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _12955_ (.A1(_04956_),
    .A2(_04959_),
    .B(_04960_),
    .ZN(_04961_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12956_ (.A1(_04208_),
    .A2(_04766_),
    .ZN(_04962_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _12957_ (.A1(_04769_),
    .A2(_04962_),
    .A3(_04763_),
    .Z(_04963_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _12958_ (.I(_04963_),
    .ZN(_04964_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12959_ (.A1(_04512_),
    .A2(_04420_),
    .ZN(_04965_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12960_ (.I(_04505_),
    .Z(_04966_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12961_ (.A1(_04486_),
    .A2(_04492_),
    .Z(_04967_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _12962_ (.A1(_04486_),
    .A2(_04492_),
    .Z(_04968_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _12963_ (.A1(_04484_),
    .A2(_04967_),
    .B(_04968_),
    .ZN(_04969_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _12964_ (.A1(_04619_),
    .A2(_04966_),
    .B(_04969_),
    .ZN(_04970_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _12965_ (.A1(_04619_),
    .A2(_04966_),
    .A3(_04969_),
    .ZN(_04971_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _12966_ (.A1(_04965_),
    .A2(_04970_),
    .B(_04971_),
    .ZN(_04972_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12967_ (.A1(_04964_),
    .A2(_04961_),
    .Z(_04973_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12968_ (.A1(_04972_),
    .A2(_04973_),
    .ZN(_04974_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _12969_ (.A1(_04961_),
    .A2(_04964_),
    .B(_04974_),
    .ZN(_04975_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12970_ (.A1(_04448_),
    .A2(_04461_),
    .ZN(_04976_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12971_ (.A1(_04808_),
    .A2(_04809_),
    .Z(_04977_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12972_ (.A1(_04976_),
    .A2(_04977_),
    .Z(_04978_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _12973_ (.A1(_04957_),
    .A2(_04956_),
    .A3(_04958_),
    .Z(_04979_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12974_ (.A1(_04976_),
    .A2(_04977_),
    .Z(_04980_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _12975_ (.A1(_04978_),
    .A2(_04979_),
    .B(_04980_),
    .ZN(_04981_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12976_ (.A1(_04811_),
    .A2(_04812_),
    .Z(_04982_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12977_ (.A1(_04981_),
    .A2(_04982_),
    .Z(_04983_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _12978_ (.A1(_04972_),
    .A2(_04973_),
    .ZN(_04984_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12979_ (.A1(_04978_),
    .A2(_04979_),
    .Z(_04985_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12980_ (.A1(_04980_),
    .A2(_04985_),
    .B(_04982_),
    .ZN(_04986_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12981_ (.A1(_04983_),
    .A2(_04984_),
    .B(_04986_),
    .ZN(_04987_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _12982_ (.A1(_04814_),
    .A2(_04870_),
    .A3(_04872_),
    .ZN(_04988_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _12983_ (.A1(_04987_),
    .A2(_04988_),
    .Z(_04989_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12984_ (.A1(_04987_),
    .A2(net52),
    .Z(_04990_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _12985_ (.A1(_04975_),
    .A2(_04989_),
    .B(_04990_),
    .ZN(_04991_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _12986_ (.A1(_04952_),
    .A2(_04991_),
    .ZN(_04992_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _12987_ (.A1(_04975_),
    .A2(_04989_),
    .ZN(_04993_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _12988_ (.A1(_04512_),
    .A2(_04642_),
    .A3(_04509_),
    .Z(_04994_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12989_ (.A1(_04503_),
    .A2(_04514_),
    .ZN(_04995_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _12990_ (.A1(_04994_),
    .A2(_04995_),
    .ZN(_04996_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12991_ (.A1(_04466_),
    .A2(_04494_),
    .Z(_04997_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _12992_ (.A1(_04465_),
    .A2(_04495_),
    .B(_04997_),
    .ZN(_04998_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12993_ (.A1(_04211_),
    .A2(_04966_),
    .ZN(_04999_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _12994_ (.A1(_04969_),
    .A2(_04999_),
    .A3(_04965_),
    .Z(_05000_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12995_ (.A1(_04998_),
    .A2(_05000_),
    .Z(_05001_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _12996_ (.I(_04998_),
    .ZN(_05002_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12997_ (.A1(_05002_),
    .A2(_05000_),
    .ZN(_05003_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _12998_ (.A1(_04996_),
    .A2(_05001_),
    .B(_05003_),
    .ZN(_05004_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _12999_ (.I(_05004_),
    .ZN(_05005_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13000_ (.A1(_04465_),
    .A2(_04495_),
    .Z(_05006_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _13001_ (.A1(_04979_),
    .A2(_04978_),
    .Z(_05007_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _13002_ (.A1(_04462_),
    .A2(_05006_),
    .B(_05007_),
    .ZN(_05008_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13003_ (.A1(_04996_),
    .A2(_05001_),
    .ZN(_05009_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13004_ (.A1(_04462_),
    .A2(_05006_),
    .A3(_05007_),
    .ZN(_05010_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _13005_ (.A1(_05008_),
    .A2(_05009_),
    .B(_05010_),
    .ZN(_05011_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _13006_ (.A1(_04984_),
    .A2(_04983_),
    .Z(_05012_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13007_ (.A1(_05011_),
    .A2(_05012_),
    .ZN(_05013_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _13008_ (.A1(_05011_),
    .A2(_05012_),
    .ZN(_05014_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13009_ (.A1(_05005_),
    .A2(_05013_),
    .B(_05014_),
    .ZN(_05015_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _13010_ (.A1(_04993_),
    .A2(_05015_),
    .Z(_05016_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _13011_ (.A1(_05011_),
    .A2(_05012_),
    .A3(_05004_),
    .ZN(_05017_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13012_ (.I(_04497_),
    .ZN(_05018_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13013_ (.A1(_04497_),
    .A2(_04515_),
    .Z(_05019_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13014_ (.A1(_04502_),
    .A2(_05019_),
    .ZN(_05020_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _13015_ (.A1(_05018_),
    .A2(_04515_),
    .B(_05020_),
    .ZN(_05021_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13016_ (.A1(_04381_),
    .A2(_04439_),
    .B(_04496_),
    .ZN(_05022_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _13017_ (.A1(_04381_),
    .A2(_04439_),
    .A3(_04496_),
    .ZN(_05023_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _13018_ (.A1(_05022_),
    .A2(_04516_),
    .B(_05023_),
    .ZN(_05024_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13019_ (.A1(_04462_),
    .A2(_05006_),
    .ZN(_05025_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _13020_ (.A1(_04996_),
    .A2(_04998_),
    .A3(_05000_),
    .Z(_05026_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _13021_ (.A1(_05025_),
    .A2(_05007_),
    .A3(_05026_),
    .Z(_05027_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13022_ (.A1(_05024_),
    .A2(_05027_),
    .ZN(_05028_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _13023_ (.A1(_05024_),
    .A2(_05027_),
    .Z(_05029_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13024_ (.A1(_05021_),
    .A2(_05028_),
    .B(_05029_),
    .ZN(_05030_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13025_ (.A1(_05017_),
    .A2(_05030_),
    .ZN(_05031_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13026_ (.A1(_05028_),
    .A2(_05021_),
    .Z(_05032_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _13027_ (.A1(_04438_),
    .A2(_04517_),
    .Z(_05033_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13028_ (.A1(_04435_),
    .A2(_04518_),
    .B(_05033_),
    .ZN(_05034_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _13029_ (.A1(_05032_),
    .A2(_05034_),
    .Z(_05035_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _13030_ (.A1(_05035_),
    .A2(_05031_),
    .ZN(_05036_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _13031_ (.A1(_04693_),
    .A2(_04992_),
    .A3(_05016_),
    .A4(_05036_),
    .ZN(_05037_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _13032_ (.A1(_05021_),
    .A2(_05028_),
    .Z(_05038_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _13033_ (.A1(_05029_),
    .A2(_05038_),
    .B(_05017_),
    .ZN(_05039_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13034_ (.A1(_05032_),
    .A2(_05034_),
    .Z(_05040_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13035_ (.A1(_05017_),
    .A2(_05029_),
    .A3(_05038_),
    .ZN(_05041_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _13036_ (.A1(_05039_),
    .A2(_05040_),
    .B(_05041_),
    .ZN(_05042_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _13037_ (.A1(_04992_),
    .A2(_05016_),
    .A3(_05042_),
    .ZN(_05043_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13038_ (.A1(_04952_),
    .A2(_04991_),
    .ZN(_05044_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _13039_ (.A1(_05011_),
    .A2(_05012_),
    .Z(_05045_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _13040_ (.A1(_05014_),
    .A2(_05004_),
    .A3(_05045_),
    .ZN(_05046_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _13041_ (.A1(_04952_),
    .A2(_04991_),
    .B1(_05014_),
    .B2(_05046_),
    .C(_04993_),
    .ZN(_05047_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _13042_ (.A1(_05044_),
    .A2(_05047_),
    .Z(_05048_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _13043_ (.I(_04923_),
    .Z(_05049_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13044_ (.A1(_04928_),
    .A2(_04930_),
    .Z(_05050_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _13045_ (.A1(_04928_),
    .A2(_04930_),
    .Z(_05051_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13046_ (.A1(_04925_),
    .A2(_05050_),
    .B(_05051_),
    .ZN(_05052_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13047_ (.A1(_04643_),
    .A2(_05049_),
    .A3(_05052_),
    .ZN(_05053_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13048_ (.I(_04946_),
    .Z(_05054_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13049_ (.A1(_04641_),
    .A2(_05049_),
    .ZN(_05055_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13050_ (.A1(_05052_),
    .A2(_05055_),
    .ZN(_05056_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13051_ (.A1(_04629_),
    .A2(_05054_),
    .A3(_05056_),
    .ZN(_05057_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13052_ (.A1(_05053_),
    .A2(_05057_),
    .Z(_05058_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _13053_ (.A1(_04917_),
    .A2(_04921_),
    .Z(_05059_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13054_ (.A1(_04922_),
    .A2(_04931_),
    .B(_05059_),
    .ZN(_05060_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13055_ (.A1(_04900_),
    .A2(_04905_),
    .ZN(_05061_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13056_ (.A1(_04900_),
    .A2(_04905_),
    .ZN(_05062_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _13057_ (.A1(_04895_),
    .A2(_05061_),
    .B(_05062_),
    .ZN(_05063_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _13058_ (.A1(_04699_),
    .A2(_04291_),
    .B1(_04511_),
    .B2(_04697_),
    .ZN(_05064_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _13059_ (.A1(_04699_),
    .A2(_04221_),
    .A3(_04274_),
    .A4(_04511_),
    .ZN(_05065_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _13060_ (.A1(_04918_),
    .A2(_05064_),
    .B(_05065_),
    .ZN(_05066_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13061_ (.A1(_04705_),
    .A2(_04751_),
    .ZN(_05067_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _13062_ (.A1(_03398_),
    .A2(_04219_),
    .A3(_04403_),
    .ZN(_05068_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _13063_ (.I(net57),
    .Z(_05069_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _13064_ (.A1(_03382_),
    .A2(_05069_),
    .A3(_04341_),
    .ZN(_05070_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13065_ (.A1(_05068_),
    .A2(_05070_),
    .ZN(_05071_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13066_ (.A1(_05071_),
    .A2(_05067_),
    .Z(_05072_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13067_ (.A1(_05066_),
    .A2(_05072_),
    .ZN(_05073_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13068_ (.I(_04926_),
    .Z(_05074_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _13069_ (.I(_05074_),
    .Z(_05075_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13070_ (.A1(_04175_),
    .A2(_05075_),
    .ZN(_05076_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13071_ (.I0(\filters.high[16] ),
    .I1(\filters.band[16] ),
    .S(_03185_),
    .Z(_05077_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13072_ (.I(_05077_),
    .Z(_05078_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _13073_ (.I(_05078_),
    .Z(_05079_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _13074_ (.A1(_04401_),
    .A2(_05079_),
    .ZN(_05080_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13075_ (.A1(_04201_),
    .A2(_04758_),
    .ZN(_05081_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _13076_ (.A1(_05076_),
    .A2(_05080_),
    .A3(_05081_),
    .Z(_05082_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13077_ (.A1(_05073_),
    .A2(_05082_),
    .ZN(_05083_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13078_ (.A1(_05063_),
    .A2(_05083_),
    .ZN(_05084_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13079_ (.A1(_05063_),
    .A2(_05083_),
    .ZN(_05085_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _13080_ (.A1(net41),
    .A2(_05084_),
    .B(_05085_),
    .ZN(_05086_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13081_ (.A1(_04288_),
    .A2(_05049_),
    .ZN(_05087_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13082_ (.A1(_05080_),
    .A2(_05081_),
    .Z(_05088_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _13083_ (.A1(_05080_),
    .A2(_05081_),
    .Z(_05089_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _13084_ (.A1(_05076_),
    .A2(_05088_),
    .B(_05089_),
    .ZN(_05090_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13085_ (.I(_04927_),
    .Z(_05091_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _13086_ (.I(_05091_),
    .Z(_05092_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13087_ (.A1(_04764_),
    .A2(_05092_),
    .ZN(_05093_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _13088_ (.A1(_05087_),
    .A2(_05090_),
    .A3(_05093_),
    .Z(_05094_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13089_ (.I(_05094_),
    .ZN(_05095_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13090_ (.A1(_05086_),
    .A2(_05095_),
    .Z(_05096_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _13091_ (.A1(_05086_),
    .A2(_05095_),
    .Z(_05097_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _13092_ (.A1(_05058_),
    .A2(_05096_),
    .B(_05097_),
    .ZN(_05098_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13093_ (.A1(_04878_),
    .A2(_04891_),
    .ZN(_05099_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13094_ (.A1(_04878_),
    .A2(_04891_),
    .ZN(_05100_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13095_ (.A1(_05099_),
    .A2(_04906_),
    .B(_05100_),
    .ZN(_05101_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13096_ (.A1(_04886_),
    .A2(_04890_),
    .ZN(_05102_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _13097_ (.A1(_04883_),
    .A2(_04885_),
    .ZN(_05103_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _13098_ (.A1(_03270_),
    .A2(_04240_),
    .A3(_04816_),
    .Z(_05104_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13099_ (.A1(_03252_),
    .A2(_04224_),
    .A3(_04880_),
    .ZN(_05105_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13100_ (.A1(\filters.cutoff_lut[16] ),
    .A2(_04441_),
    .Z(_05106_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13101_ (.I(_05106_),
    .Z(_05107_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _13102_ (.A1(_03199_),
    .A2(_04215_),
    .A3(_05107_),
    .ZN(_05108_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _13103_ (.A1(_05104_),
    .A2(_05105_),
    .A3(_05108_),
    .Z(_05109_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _13104_ (.A1(_03315_),
    .A2(_04163_),
    .A3(_04443_),
    .Z(_05110_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13105_ (.A1(net64),
    .A2(_04196_),
    .A3(_04779_),
    .ZN(_05111_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13106_ (.A1(_03301_),
    .A2(_04332_),
    .A3(_04783_),
    .ZN(_05112_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _13107_ (.A1(_05110_),
    .A2(_05111_),
    .A3(_05112_),
    .Z(_05113_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _13108_ (.A1(_05103_),
    .A2(_05109_),
    .A3(_05113_),
    .Z(_05114_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13109_ (.A1(_05102_),
    .A2(_05114_),
    .ZN(_05115_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _13110_ (.A1(_04902_),
    .A2(_04903_),
    .Z(_05116_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _13111_ (.A1(_04901_),
    .A2(_04904_),
    .B(_05116_),
    .ZN(_05117_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _13112_ (.A1(_04535_),
    .A2(_04896_),
    .ZN(_05118_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13113_ (.A1(_04888_),
    .A2(_04889_),
    .ZN(_05119_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13114_ (.A1(_04888_),
    .A2(_04889_),
    .ZN(_05120_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _13115_ (.A1(_05118_),
    .A2(_05119_),
    .B(_05120_),
    .ZN(_05121_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13116_ (.A1(_04367_),
    .A2(_04290_),
    .ZN(_05122_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13117_ (.A1(_03349_),
    .A2(_04315_),
    .A3(_04191_),
    .ZN(_05123_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _13118_ (.A1(_03332_),
    .A2(net60),
    .A3(_04450_),
    .ZN(_05124_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13119_ (.A1(_05123_),
    .A2(_05124_),
    .ZN(_05125_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13120_ (.A1(_05122_),
    .A2(_05125_),
    .ZN(_05126_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _13121_ (.A1(_05117_),
    .A2(_05121_),
    .A3(_05126_),
    .ZN(_05127_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _13122_ (.A1(_05115_),
    .A2(_05127_),
    .Z(_05128_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13123_ (.A1(_05101_),
    .A2(_05128_),
    .ZN(_05129_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _13124_ (.A1(_05060_),
    .A2(_05063_),
    .A3(_05083_),
    .ZN(_05130_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13125_ (.A1(_05101_),
    .A2(_05128_),
    .ZN(_05131_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13126_ (.A1(_05129_),
    .A2(_05130_),
    .B(_05131_),
    .ZN(_05132_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13127_ (.A1(_05102_),
    .A2(_05114_),
    .ZN(_05133_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13128_ (.A1(_05115_),
    .A2(_05127_),
    .B(_05133_),
    .ZN(_05134_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _13129_ (.A1(_05103_),
    .A2(_05109_),
    .ZN(_05135_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13130_ (.I(_05113_),
    .ZN(_05136_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13131_ (.A1(_05103_),
    .A2(_05109_),
    .ZN(_05137_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _13132_ (.A1(_05135_),
    .A2(_05136_),
    .B(_05137_),
    .ZN(_05138_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13133_ (.A1(_04369_),
    .A2(_04818_),
    .ZN(_05139_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13134_ (.A1(_05105_),
    .A2(_05108_),
    .Z(_05140_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _13135_ (.A1(_05105_),
    .A2(_05108_),
    .Z(_05141_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _13136_ (.A1(_05139_),
    .A2(_05140_),
    .B(_05141_),
    .ZN(_05142_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _13137_ (.A1(_04389_),
    .A2(_04817_),
    .ZN(_05143_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13138_ (.A1(_04368_),
    .A2(_04881_),
    .ZN(_05144_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _13139_ (.I(_05107_),
    .Z(_05145_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13140_ (.A1(_04320_),
    .A2(_05145_),
    .ZN(_05146_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _13141_ (.A1(_05143_),
    .A2(_05144_),
    .A3(_05146_),
    .ZN(_05147_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _13142_ (.A1(_04179_),
    .A2(_04800_),
    .ZN(_05148_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13143_ (.A1(_04278_),
    .A2(_04780_),
    .ZN(_05149_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13144_ (.A1(_04386_),
    .A2(_04791_),
    .ZN(_05150_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _13145_ (.A1(_05148_),
    .A2(_05149_),
    .A3(_05150_),
    .ZN(_05151_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _13146_ (.A1(_05142_),
    .A2(_05147_),
    .A3(net49),
    .Z(_05152_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _13147_ (.A1(_05123_),
    .A2(_05124_),
    .Z(_05153_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13148_ (.A1(_05122_),
    .A2(_05125_),
    .B(_05153_),
    .ZN(_05154_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13149_ (.A1(_05111_),
    .A2(_05112_),
    .Z(_05155_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _13150_ (.A1(_05111_),
    .A2(_05112_),
    .Z(_05156_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_4 _13151_ (.A1(_04165_),
    .A2(_04896_),
    .A3(_05155_),
    .B(_05156_),
    .ZN(_05157_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13152_ (.I(_04366_),
    .Z(_05158_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13153_ (.A1(_05158_),
    .A2(_04510_),
    .ZN(_05159_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13154_ (.A1(_03348_),
    .A2(_04191_),
    .A3(_04375_),
    .ZN(_05160_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13155_ (.A1(_03363_),
    .A2(_04315_),
    .A3(_04271_),
    .ZN(_05161_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13156_ (.A1(_05160_),
    .A2(_05161_),
    .ZN(_05162_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _13157_ (.A1(_05159_),
    .A2(_05162_),
    .Z(_05163_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _13158_ (.A1(_05154_),
    .A2(_05157_),
    .A3(_05163_),
    .Z(_05164_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _13159_ (.A1(_05138_),
    .A2(_05152_),
    .A3(_05164_),
    .Z(_05165_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13160_ (.A1(_05134_),
    .A2(_05165_),
    .ZN(_05166_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13161_ (.A1(_05066_),
    .A2(_05072_),
    .ZN(_05167_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _13162_ (.A1(_05073_),
    .A2(_05082_),
    .B(_05167_),
    .ZN(_05168_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13163_ (.A1(_05121_),
    .A2(_05126_),
    .ZN(_05169_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13164_ (.A1(_05121_),
    .A2(_05126_),
    .ZN(_05170_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _13165_ (.A1(_05117_),
    .A2(_05169_),
    .B(_05170_),
    .ZN(_05171_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _13166_ (.A1(_05068_),
    .A2(_05070_),
    .Z(_05172_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13167_ (.A1(_05067_),
    .A2(_05071_),
    .B(_05172_),
    .ZN(_05173_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13168_ (.A1(_04228_),
    .A2(_04737_),
    .ZN(_05174_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13169_ (.A1(_05069_),
    .A2(_04404_),
    .ZN(_05175_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13170_ (.A1(_04703_),
    .A2(_04490_),
    .ZN(_05176_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _13171_ (.A1(_05174_),
    .A2(_05175_),
    .A3(_05176_),
    .Z(_05177_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13172_ (.A1(_05173_),
    .A2(_05177_),
    .ZN(_05178_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _13173_ (.I(_03186_),
    .Z(_05179_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13174_ (.A1(\filters.band[16] ),
    .A2(_05179_),
    .Z(_05180_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _13175_ (.A1(\filters.high[16] ),
    .A2(_03470_),
    .B(_05180_),
    .ZN(_05181_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _13176_ (.A1(_05181_),
    .A2(_04537_),
    .ZN(_05182_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13177_ (.I(_04858_),
    .Z(_05183_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _13178_ (.A1(_04742_),
    .A2(_05183_),
    .ZN(_05184_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13179_ (.I0(\filters.high[17] ),
    .I1(\filters.band[17] ),
    .S(_03186_),
    .Z(_05185_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13180_ (.I(_05185_),
    .Z(_05186_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _13181_ (.I(_05186_),
    .Z(_05187_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _13182_ (.A1(_04401_),
    .A2(_05187_),
    .ZN(_05188_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _13183_ (.A1(_05182_),
    .A2(_05184_),
    .A3(_05188_),
    .Z(_05189_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13184_ (.A1(_05178_),
    .A2(_05189_),
    .ZN(_05190_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _13185_ (.A1(_05168_),
    .A2(_05171_),
    .A3(_05190_),
    .ZN(_05191_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _13186_ (.A1(_05166_),
    .A2(_05191_),
    .Z(_05192_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13187_ (.A1(_05132_),
    .A2(_05192_),
    .ZN(_05193_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _13188_ (.A1(_05058_),
    .A2(_05086_),
    .A3(_05095_),
    .Z(_05194_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13189_ (.A1(_05132_),
    .A2(_05192_),
    .ZN(_05195_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13190_ (.A1(_05193_),
    .A2(_05194_),
    .B(_05195_),
    .ZN(_05196_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13191_ (.A1(_05134_),
    .A2(_05165_),
    .ZN(_05197_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13192_ (.A1(_05166_),
    .A2(_05191_),
    .B(_05197_),
    .ZN(_05198_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13193_ (.A1(_05138_),
    .A2(_05152_),
    .ZN(_05199_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13194_ (.I(_05154_),
    .ZN(_05200_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _13195_ (.A1(_05200_),
    .A2(_05157_),
    .A3(_05163_),
    .Z(_05201_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13196_ (.A1(_05138_),
    .A2(_05152_),
    .ZN(_05202_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _13197_ (.A1(_05199_),
    .A2(_05201_),
    .B(_05202_),
    .ZN(_05203_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13198_ (.A1(_05142_),
    .A2(_05147_),
    .ZN(_05204_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13199_ (.I(_05151_),
    .ZN(_05205_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13200_ (.A1(_05142_),
    .A2(_05147_),
    .ZN(_05206_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13201_ (.A1(_05204_),
    .A2(_05205_),
    .B(_05206_),
    .ZN(_05207_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _13202_ (.I(_05107_),
    .Z(_05208_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _13203_ (.A1(_04369_),
    .A2(_04882_),
    .B1(_05208_),
    .B2(_04320_),
    .ZN(_05209_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _13204_ (.A1(_04320_),
    .A2(_04368_),
    .A3(_04882_),
    .A4(_05145_),
    .ZN(_05210_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _13205_ (.A1(_05143_),
    .A2(_05209_),
    .B(_05210_),
    .ZN(_05211_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13206_ (.A1(_04277_),
    .A2(_04817_),
    .ZN(_05212_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13207_ (.A1(_03285_),
    .A2(_04195_),
    .A3(_04880_),
    .ZN(_05213_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13208_ (.A1(_03270_),
    .A2(_04240_),
    .A3(_05106_),
    .ZN(_05214_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13209_ (.A1(_05213_),
    .A2(_05214_),
    .ZN(_05215_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _13210_ (.A1(_05212_),
    .A2(_05215_),
    .Z(_05216_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13211_ (.A1(_05211_),
    .A2(_05216_),
    .ZN(_05217_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13212_ (.A1(_04485_),
    .A2(_04444_),
    .ZN(_05218_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _13213_ (.A1(_04386_),
    .A2(_04180_),
    .A3(_04824_),
    .A4(_04791_),
    .Z(_05219_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _13214_ (.I(_04780_),
    .Z(_05220_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _13215_ (.A1(_04386_),
    .A2(_05220_),
    .B1(_04791_),
    .B2(_04180_),
    .ZN(_05221_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _13216_ (.A1(_05218_),
    .A2(_05219_),
    .A3(_05221_),
    .Z(_05222_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13217_ (.A1(_05219_),
    .A2(_05221_),
    .B(_05218_),
    .ZN(_05223_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _13218_ (.A1(_05222_),
    .A2(_05223_),
    .ZN(_05224_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _13219_ (.A1(_05224_),
    .A2(_05217_),
    .Z(_05225_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13220_ (.A1(_05160_),
    .A2(_05161_),
    .ZN(_05226_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13221_ (.A1(_05159_),
    .A2(_05162_),
    .ZN(_05227_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13222_ (.A1(_05227_),
    .A2(_05226_),
    .ZN(_05228_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13223_ (.I(_04824_),
    .Z(_05229_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _13224_ (.I(_04784_),
    .Z(_05230_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _13225_ (.I(_04385_),
    .Z(_05231_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _13226_ (.A1(_04280_),
    .A2(_05229_),
    .B1(_05230_),
    .B2(_05231_),
    .ZN(_05232_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _13227_ (.A1(_04280_),
    .A2(_05231_),
    .A3(_04825_),
    .A4(_05230_),
    .ZN(_05233_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _13228_ (.A1(_05148_),
    .A2(_05232_),
    .B(_05233_),
    .ZN(_05234_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13229_ (.A1(_04324_),
    .A2(_04405_),
    .Z(_05235_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _13230_ (.A1(_03363_),
    .A2(_04271_),
    .A3(_04450_),
    .ZN(_05236_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _13231_ (.A1(_03382_),
    .A2(_04371_),
    .A3(_04342_),
    .ZN(_05237_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13232_ (.A1(_05236_),
    .A2(_05237_),
    .Z(_05238_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13233_ (.A1(_05235_),
    .A2(_05238_),
    .Z(_05239_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _13234_ (.A1(_05228_),
    .A2(_05234_),
    .A3(_05239_),
    .ZN(_05240_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _13235_ (.A1(_05207_),
    .A2(_05225_),
    .A3(_05240_),
    .Z(_05241_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _13236_ (.A1(_05067_),
    .A2(_05071_),
    .Z(_05242_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _13237_ (.A1(_05172_),
    .A2(_05242_),
    .B(_05177_),
    .ZN(_05243_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _13238_ (.A1(_05178_),
    .A2(_05189_),
    .B(_05243_),
    .ZN(_05244_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13239_ (.A1(_05157_),
    .A2(_05163_),
    .ZN(_05245_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13240_ (.A1(_05157_),
    .A2(_05163_),
    .ZN(_05246_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13241_ (.A1(_05200_),
    .A2(_05245_),
    .B(_05246_),
    .ZN(_05247_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _13242_ (.A1(_04255_),
    .A2(_04864_),
    .B1(_04491_),
    .B2(_04471_),
    .ZN(_05248_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _13243_ (.A1(_04255_),
    .A2(_04392_),
    .A3(_04405_),
    .A4(_04751_),
    .ZN(_05249_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _13244_ (.A1(_05174_),
    .A2(_05248_),
    .B(_05249_),
    .ZN(_05250_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13245_ (.A1(_04228_),
    .A2(_04740_),
    .ZN(_05251_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13246_ (.A1(_05069_),
    .A2(_04750_),
    .ZN(_05252_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13247_ (.A1(_04470_),
    .A2(_04712_),
    .ZN(_05253_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _13248_ (.A1(_05251_),
    .A2(_05252_),
    .A3(_05253_),
    .Z(_05254_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13249_ (.A1(_05250_),
    .A2(_05254_),
    .ZN(_05255_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13250_ (.I(_05186_),
    .Z(_05256_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13251_ (.A1(_04266_),
    .A2(_05256_),
    .ZN(_05257_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13252_ (.A1(_04199_),
    .A2(_04862_),
    .ZN(_05258_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13253_ (.I0(\filters.high[18] ),
    .I1(\filters.band[18] ),
    .S(_03185_),
    .Z(_05259_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13254_ (.I(_05259_),
    .Z(_05260_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13255_ (.A1(_04185_),
    .A2(_05260_),
    .ZN(_05261_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13256_ (.A1(_05258_),
    .A2(_05261_),
    .Z(_05262_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _13257_ (.A1(_05257_),
    .A2(_05262_),
    .ZN(_05263_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13258_ (.A1(_05255_),
    .A2(_05263_),
    .Z(_05264_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _13259_ (.A1(_05244_),
    .A2(_05247_),
    .A3(_05264_),
    .ZN(_05265_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _13260_ (.A1(_05203_),
    .A2(_05241_),
    .A3(_05265_),
    .Z(_05266_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13261_ (.A1(_05198_),
    .A2(_05266_),
    .ZN(_05267_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _13262_ (.I(_05092_),
    .Z(_05268_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _13263_ (.A1(_04765_),
    .A2(_05268_),
    .B(_05090_),
    .ZN(_05269_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13264_ (.A1(_04765_),
    .A2(_05268_),
    .A3(_05090_),
    .ZN(_05270_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13265_ (.A1(_05087_),
    .A2(_05269_),
    .B(_05270_),
    .ZN(_05271_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13266_ (.A1(_05171_),
    .A2(_05190_),
    .ZN(_05272_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13267_ (.A1(_05171_),
    .A2(_05190_),
    .ZN(_05273_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _13268_ (.A1(_05168_),
    .A2(_05272_),
    .B(_05273_),
    .ZN(_05274_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13269_ (.A1(_04629_),
    .A2(_05268_),
    .ZN(_05275_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13270_ (.A1(_05184_),
    .A2(_05188_),
    .ZN(_05276_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13271_ (.A1(_05184_),
    .A2(_05188_),
    .ZN(_05277_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _13272_ (.A1(net48),
    .A2(_05276_),
    .B(_05277_),
    .ZN(_05278_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13273_ (.I(_05077_),
    .Z(_05279_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13274_ (.I(_05279_),
    .Z(_05280_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _13275_ (.I(_05280_),
    .Z(_05281_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13276_ (.A1(_04302_),
    .A2(_05281_),
    .ZN(_05282_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13277_ (.A1(_05278_),
    .A2(_05282_),
    .Z(_05283_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13278_ (.A1(_05275_),
    .A2(_05283_),
    .ZN(_05284_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _13279_ (.A1(_05271_),
    .A2(_05274_),
    .A3(_05284_),
    .Z(_05285_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13280_ (.A1(_05267_),
    .A2(_05285_),
    .Z(_05286_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13281_ (.A1(_05196_),
    .A2(_05286_),
    .Z(_05287_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13282_ (.A1(_05196_),
    .A2(_05286_),
    .Z(_05288_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _13283_ (.A1(_05098_),
    .A2(net45),
    .B(_05288_),
    .ZN(_05289_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13284_ (.I(_05284_),
    .ZN(_05290_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13285_ (.A1(_05274_),
    .A2(_05290_),
    .Z(_05291_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13286_ (.A1(_05271_),
    .A2(_05291_),
    .ZN(_05292_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13287_ (.A1(_05274_),
    .A2(_05290_),
    .B(_05292_),
    .ZN(_05293_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13288_ (.A1(_05198_),
    .A2(_05266_),
    .ZN(_05294_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13289_ (.A1(_05267_),
    .A2(_05285_),
    .B(_05294_),
    .ZN(_05295_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13290_ (.A1(_05203_),
    .A2(_05241_),
    .ZN(_05296_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13291_ (.I(_05265_),
    .ZN(_05297_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13292_ (.A1(_05203_),
    .A2(_05241_),
    .ZN(_05298_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _13293_ (.A1(_05296_),
    .A2(_05297_),
    .B(_05298_),
    .ZN(_05299_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13294_ (.A1(_05207_),
    .A2(_05225_),
    .ZN(_05300_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13295_ (.I(_05240_),
    .ZN(_05301_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13296_ (.A1(_05207_),
    .A2(_05225_),
    .ZN(_05302_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13297_ (.A1(_05300_),
    .A2(_05301_),
    .B(_05302_),
    .ZN(_05303_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13298_ (.A1(_05211_),
    .A2(_05216_),
    .ZN(_05304_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13299_ (.A1(_05217_),
    .A2(_05224_),
    .B(_05304_),
    .ZN(_05305_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _13300_ (.A1(_05213_),
    .A2(_05214_),
    .Z(_05306_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13301_ (.A1(_05212_),
    .A2(_05215_),
    .B(_05306_),
    .ZN(_05307_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13302_ (.A1(_04384_),
    .A2(_04816_),
    .ZN(_05308_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13303_ (.A1(_03300_),
    .A2(_04276_),
    .A3(_04879_),
    .ZN(_05309_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13304_ (.A1(_03285_),
    .A2(_04194_),
    .A3(_05106_),
    .ZN(_05310_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13305_ (.A1(_05309_),
    .A2(_05310_),
    .ZN(_05311_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13306_ (.A1(_05308_),
    .A2(_05311_),
    .Z(_05312_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _13307_ (.A1(_05307_),
    .A2(_05312_),
    .ZN(_05313_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13308_ (.A1(_04273_),
    .A2(_04800_),
    .ZN(_05314_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _13309_ (.A1(_04267_),
    .A2(_04179_),
    .A3(_04781_),
    .A4(_04803_),
    .Z(_05315_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _13310_ (.A1(_04477_),
    .A2(_04781_),
    .B1(_04784_),
    .B2(_04267_),
    .ZN(_05316_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _13311_ (.A1(_05314_),
    .A2(_05315_),
    .A3(_05316_),
    .Z(_05317_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13312_ (.A1(_05315_),
    .A2(_05316_),
    .B(_05314_),
    .ZN(_05318_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13313_ (.A1(_05317_),
    .A2(_05318_),
    .ZN(_05319_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13314_ (.A1(_05313_),
    .A2(_05319_),
    .Z(_05320_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13315_ (.A1(_05320_),
    .A2(_05305_),
    .ZN(_05321_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13316_ (.A1(_05235_),
    .A2(_05238_),
    .ZN(_05322_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _13317_ (.A1(_05236_),
    .A2(_05237_),
    .B(_05322_),
    .ZN(_05323_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _13318_ (.A1(_04695_),
    .A2(_04729_),
    .A3(_05220_),
    .A4(_04804_),
    .ZN(_05324_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13319_ (.A1(_05218_),
    .A2(_05221_),
    .B(_05324_),
    .ZN(_05325_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13320_ (.A1(_04323_),
    .A2(_04489_),
    .ZN(_05326_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13321_ (.A1(_04395_),
    .A2(_04375_),
    .ZN(_05327_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13322_ (.A1(_04315_),
    .A2(_04404_),
    .ZN(_05328_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _13323_ (.A1(_05326_),
    .A2(_05327_),
    .A3(_05328_),
    .Z(_05329_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13324_ (.A1(_05329_),
    .A2(_05325_),
    .ZN(_05330_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13325_ (.A1(_05323_),
    .A2(_05330_),
    .ZN(_05331_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13326_ (.A1(_05331_),
    .A2(_05321_),
    .Z(_05332_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13327_ (.I(_05250_),
    .ZN(_05333_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13328_ (.A1(_05255_),
    .A2(_05263_),
    .ZN(_05334_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _13329_ (.A1(_05333_),
    .A2(_05254_),
    .B(_05334_),
    .ZN(_05335_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13330_ (.A1(_05234_),
    .A2(_05239_),
    .ZN(_05336_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13331_ (.A1(_05234_),
    .A2(_05239_),
    .ZN(_05337_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13332_ (.A1(net69),
    .A2(_05336_),
    .B(_05337_),
    .ZN(_05338_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _13333_ (.A1(net68),
    .A2(_04490_),
    .B1(_04712_),
    .B2(_04703_),
    .ZN(_05339_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _13334_ (.A1(_04254_),
    .A2(_04470_),
    .A3(_04490_),
    .A4(_04712_),
    .ZN(_05340_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _13335_ (.A1(_05251_),
    .A2(_05339_),
    .B(_05340_),
    .ZN(_05341_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13336_ (.A1(_04227_),
    .A2(_04860_),
    .ZN(_05342_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13337_ (.A1(net57),
    .A2(_04711_),
    .ZN(_05343_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13338_ (.A1(_04257_),
    .A2(_04739_),
    .ZN(_05344_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _13339_ (.A1(_05342_),
    .A2(_05343_),
    .A3(_05344_),
    .Z(_05345_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13340_ (.A1(_05341_),
    .A2(_05345_),
    .ZN(_05346_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13341_ (.I(_05259_),
    .Z(_05347_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13342_ (.A1(_04265_),
    .A2(_05347_),
    .ZN(_05348_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13343_ (.A1(_04198_),
    .A2(_04926_),
    .ZN(_05349_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13344_ (.I0(\filters.high[19] ),
    .I1(\filters.band[19] ),
    .S(_04710_),
    .Z(_05350_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13345_ (.I(_05350_),
    .Z(_05351_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13346_ (.A1(_04184_),
    .A2(_05351_),
    .ZN(_05352_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13347_ (.A1(_05349_),
    .A2(_05352_),
    .Z(_05353_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _13348_ (.A1(_05348_),
    .A2(_05353_),
    .ZN(_05354_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13349_ (.A1(_05346_),
    .A2(_05354_),
    .Z(_05355_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13350_ (.A1(_05338_),
    .A2(_05355_),
    .Z(_05356_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _13351_ (.A1(_05335_),
    .A2(_05356_),
    .Z(_05357_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _13352_ (.A1(_05303_),
    .A2(_05332_),
    .A3(_05357_),
    .Z(_05358_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13353_ (.A1(_04500_),
    .A2(_05092_),
    .A3(_05283_),
    .ZN(_05359_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _13354_ (.A1(_05278_),
    .A2(_05282_),
    .B(_05359_),
    .ZN(_05360_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13355_ (.I(_05244_),
    .ZN(_05361_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _13356_ (.A1(_05247_),
    .A2(_05264_),
    .Z(_05362_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13357_ (.A1(_05247_),
    .A2(_05264_),
    .Z(_05363_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _13358_ (.A1(_05361_),
    .A2(_05362_),
    .B(_05363_),
    .ZN(_05364_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13359_ (.A1(_04420_),
    .A2(_05281_),
    .ZN(_05365_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _13360_ (.A1(_05258_),
    .A2(_05261_),
    .Z(_05366_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13361_ (.I(_05187_),
    .Z(_05367_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13362_ (.A1(_04596_),
    .A2(_05367_),
    .A3(_05262_),
    .ZN(_05368_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13363_ (.A1(_05366_),
    .A2(_05368_),
    .Z(_05369_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13364_ (.I(_05367_),
    .Z(_05370_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13365_ (.A1(_04641_),
    .A2(_05370_),
    .ZN(_05371_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _13366_ (.A1(_05369_),
    .A2(_05371_),
    .Z(_05372_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13367_ (.A1(_05365_),
    .A2(_05372_),
    .Z(_05373_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _13368_ (.A1(_05360_),
    .A2(_05364_),
    .A3(_05373_),
    .Z(_05374_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _13369_ (.A1(_05299_),
    .A2(_05358_),
    .A3(_05374_),
    .ZN(_05375_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13370_ (.A1(_05375_),
    .A2(_05295_),
    .ZN(_05376_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _13371_ (.A1(_05376_),
    .A2(_05293_),
    .ZN(_05377_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13372_ (.A1(_05289_),
    .A2(_05377_),
    .ZN(_05378_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _13373_ (.A1(_05098_),
    .A2(_05287_),
    .ZN(_05379_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13374_ (.A1(_04914_),
    .A2(_04932_),
    .ZN(_05380_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13375_ (.A1(_04914_),
    .A2(_04932_),
    .ZN(_05381_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _13376_ (.A1(_04911_),
    .A2(_05380_),
    .B(_05381_),
    .ZN(_05382_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13377_ (.A1(_04629_),
    .A2(_05054_),
    .ZN(_05383_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13378_ (.A1(_05383_),
    .A2(_05056_),
    .ZN(_05384_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13379_ (.I(_05384_),
    .ZN(_05385_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _13380_ (.A1(_04643_),
    .A2(_05054_),
    .B(_04944_),
    .ZN(_05386_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13381_ (.A1(_04643_),
    .A2(_05054_),
    .A3(_04944_),
    .ZN(_05387_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13382_ (.A1(_04941_),
    .A2(_05386_),
    .B(_05387_),
    .ZN(_05388_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13383_ (.A1(_05382_),
    .A2(_05385_),
    .Z(_05389_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13384_ (.A1(_05388_),
    .A2(_05389_),
    .ZN(_05390_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _13385_ (.A1(_05382_),
    .A2(_05385_),
    .B(_05390_),
    .ZN(_05391_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13386_ (.A1(_04877_),
    .A2(_04907_),
    .ZN(_05392_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13387_ (.A1(_04877_),
    .A2(_04907_),
    .ZN(_05393_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _13388_ (.A1(_05392_),
    .A2(_04933_),
    .B(_05393_),
    .ZN(_05394_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _13389_ (.A1(_05129_),
    .A2(_05130_),
    .Z(_05395_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13390_ (.A1(_05394_),
    .A2(_05395_),
    .ZN(_05396_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _13391_ (.A1(_05388_),
    .A2(_05382_),
    .A3(_05384_),
    .Z(_05397_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13392_ (.A1(_05394_),
    .A2(_05395_),
    .ZN(_05398_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13393_ (.A1(_05396_),
    .A2(_05397_),
    .B(_05398_),
    .ZN(_05399_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _13394_ (.A1(_05132_),
    .A2(_05192_),
    .A3(_05194_),
    .ZN(_05400_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _13395_ (.A1(_05399_),
    .A2(_05400_),
    .Z(_05401_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13396_ (.A1(_05399_),
    .A2(_05400_),
    .Z(_05402_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _13397_ (.A1(_05391_),
    .A2(_05401_),
    .B(_05402_),
    .ZN(_05403_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _13398_ (.A1(_05403_),
    .A2(_05379_),
    .ZN(_05404_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _13399_ (.A1(_05391_),
    .A2(_05401_),
    .ZN(_05405_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13400_ (.I(_04940_),
    .ZN(_05406_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13401_ (.A1(_05406_),
    .A2(_04948_),
    .ZN(_05407_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13402_ (.A1(_04938_),
    .A2(_04949_),
    .ZN(_05408_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _13403_ (.A1(_05407_),
    .A2(_05408_),
    .ZN(_05409_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _13404_ (.A1(_04876_),
    .A2(_04934_),
    .Z(_05410_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13405_ (.A1(_04935_),
    .A2(_04950_),
    .B(_05410_),
    .ZN(_05411_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _13406_ (.A1(_05394_),
    .A2(_05395_),
    .A3(_05397_),
    .ZN(_05412_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _13407_ (.A1(_05412_),
    .A2(_05411_),
    .Z(_05413_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13408_ (.A1(net61),
    .A2(_05412_),
    .Z(_05414_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _13409_ (.A1(_05409_),
    .A2(net66),
    .B(_05414_),
    .ZN(_05415_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _13410_ (.A1(_05405_),
    .A2(_05415_),
    .ZN(_05416_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _13411_ (.A1(_05413_),
    .A2(_05409_),
    .ZN(_05417_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _13412_ (.A1(_04874_),
    .A2(_04951_),
    .Z(_05418_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13413_ (.A1(_04874_),
    .A2(_04951_),
    .Z(_05419_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _13414_ (.A1(_04775_),
    .A2(_05418_),
    .B(_05419_),
    .ZN(_05420_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _13415_ (.A1(_05417_),
    .A2(_05420_),
    .ZN(_05421_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _13416_ (.A1(net55),
    .A2(_05404_),
    .A3(_05416_),
    .A4(_05421_),
    .ZN(_05422_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_4 _13417_ (.A1(_05037_),
    .A2(_05043_),
    .A3(_05048_),
    .B(_05422_),
    .ZN(_05423_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13418_ (.A1(_05289_),
    .A2(_05377_),
    .ZN(_05424_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _13419_ (.A1(_05379_),
    .A2(_05403_),
    .ZN(_05425_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _13420_ (.A1(_05378_),
    .A2(_05404_),
    .ZN(_05426_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13421_ (.A1(_05405_),
    .A2(_05415_),
    .ZN(_05427_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _13422_ (.A1(_05405_),
    .A2(_05415_),
    .B1(_05417_),
    .B2(_05420_),
    .ZN(_05428_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13423_ (.A1(_05427_),
    .A2(_05428_),
    .Z(_05429_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13424_ (.A1(_05289_),
    .A2(_05377_),
    .ZN(_05430_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _13425_ (.A1(_05424_),
    .A2(_05425_),
    .B1(_05426_),
    .B2(_05429_),
    .C(_05430_),
    .ZN(_05431_));
 gf180mcu_fd_sc_mcu7t5v0__and2_4 _13426_ (.A1(_05423_),
    .A2(_05431_),
    .Z(_05432_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13427_ (.A1(_05364_),
    .A2(_05373_),
    .ZN(_05433_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13428_ (.A1(_05364_),
    .A2(_05373_),
    .ZN(_05434_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _13429_ (.A1(_05360_),
    .A2(_05433_),
    .B(_05434_),
    .ZN(_05435_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13430_ (.A1(_05299_),
    .A2(_05358_),
    .ZN(_05436_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13431_ (.I(_05374_),
    .ZN(_05437_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13432_ (.A1(_05299_),
    .A2(_05358_),
    .ZN(_05438_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _13433_ (.A1(_05436_),
    .A2(_05437_),
    .B(_05438_),
    .ZN(_05439_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _13434_ (.I(_04562_),
    .Z(_05440_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13435_ (.A1(_05440_),
    .A2(_05281_),
    .A3(_05372_),
    .ZN(_05441_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _13436_ (.A1(_05369_),
    .A2(_05371_),
    .B(_05441_),
    .ZN(_05442_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13437_ (.A1(_05338_),
    .A2(_05355_),
    .Z(_05443_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _13438_ (.A1(_05335_),
    .A2(_05356_),
    .B(_05443_),
    .ZN(_05444_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13439_ (.A1(_04561_),
    .A2(_05370_),
    .ZN(_05445_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _13440_ (.I(_04596_),
    .Z(_05446_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13441_ (.I(_05260_),
    .Z(_05447_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13442_ (.I(_05447_),
    .Z(_05448_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13443_ (.I(_05448_),
    .Z(_05449_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13444_ (.A1(_05446_),
    .A2(_05449_),
    .A3(_05353_),
    .ZN(_05450_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _13445_ (.A1(_05349_),
    .A2(_05352_),
    .B(_05450_),
    .ZN(_05451_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13446_ (.A1(_04642_),
    .A2(_05449_),
    .ZN(_05452_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13447_ (.A1(_05451_),
    .A2(_05452_),
    .ZN(_05453_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13448_ (.A1(_05445_),
    .A2(_05453_),
    .Z(_05454_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13449_ (.A1(_05444_),
    .A2(_05454_),
    .Z(_05455_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13450_ (.A1(_05442_),
    .A2(_05455_),
    .ZN(_05456_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _13451_ (.A1(_05303_),
    .A2(_05332_),
    .Z(_05457_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13452_ (.A1(_05303_),
    .A2(_05332_),
    .Z(_05458_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _13453_ (.A1(_05457_),
    .A2(_05357_),
    .B(_05458_),
    .ZN(_05459_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13454_ (.A1(_05305_),
    .A2(_05320_),
    .ZN(_05460_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13455_ (.A1(_05321_),
    .A2(_05331_),
    .B(_05460_),
    .ZN(_05461_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13456_ (.A1(_05327_),
    .A2(_05328_),
    .Z(_05462_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _13457_ (.A1(_05327_),
    .A2(_05328_),
    .Z(_05463_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _13458_ (.A1(_05326_),
    .A2(_05462_),
    .B(_05463_),
    .ZN(_05464_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _13459_ (.I(_05229_),
    .Z(_05465_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _13460_ (.I(_04805_),
    .Z(_05466_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _13461_ (.A1(_04269_),
    .A2(_04182_),
    .A3(_05465_),
    .A4(_05466_),
    .ZN(_05467_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13462_ (.A1(_05314_),
    .A2(_05316_),
    .B(_05467_),
    .ZN(_05468_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _13463_ (.I(_04737_),
    .Z(_05469_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13464_ (.A1(_05158_),
    .A2(_05469_),
    .ZN(_05470_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13465_ (.A1(_04451_),
    .A2(_04405_),
    .ZN(_05471_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13466_ (.A1(_04317_),
    .A2(_04752_),
    .ZN(_05472_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _13467_ (.A1(_05470_),
    .A2(_05471_),
    .A3(_05472_),
    .Z(_05473_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13468_ (.A1(_05468_),
    .A2(_05473_),
    .ZN(_05474_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13469_ (.A1(_05474_),
    .A2(_05464_),
    .ZN(_05475_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13470_ (.A1(_05307_),
    .A2(_05312_),
    .ZN(_05476_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13471_ (.A1(_05313_),
    .A2(_05319_),
    .B(_05476_),
    .ZN(_05477_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13472_ (.A1(_04511_),
    .A2(_04445_),
    .ZN(_05478_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _13473_ (.A1(_03350_),
    .A2(_04192_),
    .A3(_05220_),
    .ZN(_05479_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _13474_ (.A1(_03364_),
    .A2(_04854_),
    .A3(_04804_),
    .ZN(_05480_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13475_ (.A1(_05479_),
    .A2(_05480_),
    .Z(_05481_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13476_ (.A1(_05478_),
    .A2(_05481_),
    .Z(_05482_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _13477_ (.A1(_05309_),
    .A2(_05310_),
    .Z(_05483_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _13478_ (.A1(_05308_),
    .A2(_05311_),
    .B(_05483_),
    .ZN(_05484_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13479_ (.A1(_04477_),
    .A2(_04884_),
    .ZN(_05485_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13480_ (.A1(_04278_),
    .A2(_05208_),
    .ZN(_05486_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _13481_ (.I(_04882_),
    .Z(_05487_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13482_ (.A1(_04480_),
    .A2(_05487_),
    .ZN(_05488_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _13483_ (.A1(_05485_),
    .A2(_05486_),
    .A3(_05488_),
    .ZN(_05489_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13484_ (.A1(_05484_),
    .A2(_05489_),
    .ZN(_05490_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13485_ (.A1(_05482_),
    .A2(_05490_),
    .Z(_05491_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13486_ (.A1(_05477_),
    .A2(_05491_),
    .ZN(_05492_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13487_ (.A1(_05475_),
    .A2(_05492_),
    .Z(_05493_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _13488_ (.A1(_05461_),
    .A2(_05493_),
    .Z(_05494_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13489_ (.I(_05341_),
    .ZN(_05495_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13490_ (.A1(_05495_),
    .A2(_05345_),
    .ZN(_05496_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _13491_ (.A1(_05346_),
    .A2(_05354_),
    .B(_05496_),
    .ZN(_05497_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _13492_ (.A1(_05324_),
    .A2(_05222_),
    .B(_05329_),
    .ZN(_05498_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _13493_ (.A1(_05323_),
    .A2(net47),
    .B(_05498_),
    .ZN(_05499_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13494_ (.I(_05351_),
    .Z(_05500_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13495_ (.I(_05500_),
    .Z(_05501_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13496_ (.A1(_04525_),
    .A2(_05501_),
    .ZN(_05502_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13497_ (.A1(_04295_),
    .A2(_05279_),
    .ZN(_05503_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13498_ (.I0(\filters.high[20] ),
    .I1(\filters.band[20] ),
    .S(_03186_),
    .Z(_05504_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13499_ (.I(_05504_),
    .Z(_05505_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13500_ (.A1(_04401_),
    .A2(_05505_),
    .ZN(_05506_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13501_ (.A1(_05503_),
    .A2(_05506_),
    .Z(_05507_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13502_ (.A1(_05502_),
    .A2(_05507_),
    .ZN(_05508_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _13503_ (.I(_04848_),
    .Z(_05509_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _13504_ (.I(_04850_),
    .Z(_05510_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _13505_ (.A1(_05509_),
    .A2(_04758_),
    .B1(_04946_),
    .B2(_05510_),
    .ZN(_05511_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _13506_ (.I(_04467_),
    .Z(_05512_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _13507_ (.A1(_05512_),
    .A2(_05510_),
    .A3(_04758_),
    .A4(_04946_),
    .ZN(_05513_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _13508_ (.A1(_05342_),
    .A2(_05511_),
    .B(_05513_),
    .ZN(_05514_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13509_ (.A1(_04705_),
    .A2(_05074_),
    .ZN(_05515_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13510_ (.I(_04740_),
    .Z(_05516_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13511_ (.A1(_04237_),
    .A2(_05516_),
    .ZN(_05517_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13512_ (.I(_04862_),
    .Z(_05518_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13513_ (.A1(_04850_),
    .A2(_05518_),
    .ZN(_05519_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _13514_ (.A1(_05515_),
    .A2(_05517_),
    .A3(_05519_),
    .Z(_05520_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13515_ (.A1(_05514_),
    .A2(_05520_),
    .ZN(_05521_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13516_ (.A1(_05508_),
    .A2(_05521_),
    .ZN(_05522_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13517_ (.A1(_05499_),
    .A2(_05522_),
    .ZN(_05523_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13518_ (.A1(_05497_),
    .A2(_05523_),
    .Z(_05524_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13519_ (.A1(_05494_),
    .A2(_05524_),
    .Z(_05525_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _13520_ (.A1(_05456_),
    .A2(_05459_),
    .A3(_05525_),
    .Z(_05526_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _13521_ (.A1(_05435_),
    .A2(_05439_),
    .A3(_05526_),
    .ZN(_05527_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13522_ (.I(_05295_),
    .ZN(_05528_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13523_ (.A1(_05293_),
    .A2(_05376_),
    .ZN(_05529_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _13524_ (.A1(_05528_),
    .A2(net44),
    .B(_05529_),
    .ZN(_05530_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _13525_ (.A1(_05527_),
    .A2(_05530_),
    .ZN(_05531_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _13526_ (.A1(_05531_),
    .A2(_05432_),
    .Z(_05532_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _13527_ (.I(_05532_),
    .Z(_05533_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13528_ (.I(\filters.low[0] ),
    .Z(_05534_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13529_ (.A1(_05534_),
    .A2(_03346_),
    .ZN(_05535_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13530_ (.A1(\filters.band[0] ),
    .A2(_03471_),
    .ZN(_05536_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _13531_ (.A1(_05533_),
    .A2(_05535_),
    .A3(_05536_),
    .Z(_05537_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _13532_ (.A1(_05535_),
    .A2(_05536_),
    .B(_05533_),
    .ZN(_05538_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13533_ (.A1(_05537_),
    .A2(_05538_),
    .ZN(_05539_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13534_ (.I(_04159_),
    .Z(_05540_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13535_ (.I(_03721_),
    .Z(_05541_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13536_ (.A1(\filters.band[0] ),
    .A2(_05540_),
    .B(_05541_),
    .ZN(_05542_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _13537_ (.A1(_04161_),
    .A2(_05539_),
    .B(_05542_),
    .ZN(_00526_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _13538_ (.A1(_03730_),
    .A2(_03477_),
    .ZN(_05543_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13539_ (.I(_05543_),
    .Z(_05544_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13540_ (.I(_05544_),
    .Z(_05545_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _13541_ (.I(_05543_),
    .Z(_05546_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _13542_ (.I(_05546_),
    .Z(_05547_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13543_ (.A1(_05533_),
    .A2(_05535_),
    .A3(_05536_),
    .ZN(_05548_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13544_ (.A1(_05527_),
    .A2(_05530_),
    .Z(_05549_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _13545_ (.A1(net35),
    .A2(net39),
    .B(_05531_),
    .ZN(_05550_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13546_ (.A1(_05439_),
    .A2(_05526_),
    .ZN(_05551_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13547_ (.A1(_05439_),
    .A2(_05526_),
    .ZN(_05552_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _13548_ (.A1(_05435_),
    .A2(_05551_),
    .B(_05552_),
    .ZN(_05553_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13549_ (.A1(_05444_),
    .A2(_05454_),
    .ZN(_05554_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _13550_ (.A1(_05442_),
    .A2(_05455_),
    .B(_05554_),
    .ZN(_05555_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13551_ (.A1(_05494_),
    .A2(_05524_),
    .Z(_05556_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13552_ (.A1(_05494_),
    .A2(_05524_),
    .ZN(_05557_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13553_ (.A1(_05459_),
    .A2(_05525_),
    .Z(_05558_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _13554_ (.A1(_05459_),
    .A2(_05556_),
    .A3(_05557_),
    .B1(_05558_),
    .B2(_05456_),
    .ZN(_05559_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _13555_ (.I(_04645_),
    .Z(_05560_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13556_ (.I(_05449_),
    .Z(_05561_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13557_ (.A1(_05560_),
    .A2(_05561_),
    .A3(_05451_),
    .ZN(_05562_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _13558_ (.I(_04562_),
    .Z(_05563_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13559_ (.A1(_05563_),
    .A2(_05370_),
    .A3(_05453_),
    .ZN(_05564_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13560_ (.A1(_05562_),
    .A2(_05564_),
    .Z(_05565_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13561_ (.A1(_05499_),
    .A2(_05522_),
    .ZN(_05566_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13562_ (.A1(_05497_),
    .A2(_05523_),
    .ZN(_05567_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13563_ (.A1(_05566_),
    .A2(_05567_),
    .ZN(_05568_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13564_ (.A1(_04630_),
    .A2(_05561_),
    .ZN(_05569_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13565_ (.I(_05501_),
    .Z(_05570_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13566_ (.A1(_04597_),
    .A2(_05570_),
    .A3(_05507_),
    .ZN(_05571_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13567_ (.A1(_05503_),
    .A2(_05506_),
    .B(_05571_),
    .ZN(_05572_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13568_ (.A1(_04764_),
    .A2(_05570_),
    .ZN(_05573_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13569_ (.A1(_05572_),
    .A2(_05573_),
    .ZN(_05574_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13570_ (.A1(_05569_),
    .A2(_05574_),
    .Z(_05575_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13571_ (.A1(_05568_),
    .A2(_05575_),
    .ZN(_05576_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13572_ (.A1(_05565_),
    .A2(_05576_),
    .Z(_05577_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13573_ (.A1(_05461_),
    .A2(_05493_),
    .Z(_05578_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _13574_ (.A1(_05494_),
    .A2(_05524_),
    .B(_05578_),
    .ZN(_05579_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13575_ (.I(_05514_),
    .ZN(_05580_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13576_ (.A1(_05580_),
    .A2(_05520_),
    .ZN(_05581_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _13577_ (.A1(_05508_),
    .A2(_05521_),
    .B(_05581_),
    .ZN(_05582_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _13578_ (.A1(_05467_),
    .A2(_05317_),
    .B(_05473_),
    .ZN(_05583_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _13579_ (.A1(_05464_),
    .A2(_05474_),
    .B(_05583_),
    .ZN(_05584_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13580_ (.I(_05504_),
    .Z(_05585_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13581_ (.A1(_04176_),
    .A2(_05585_),
    .ZN(_05586_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13582_ (.A1(_04294_),
    .A2(_05186_),
    .ZN(_05587_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13583_ (.I0(\filters.high[21] ),
    .I1(\filters.band[21] ),
    .S(_05179_),
    .Z(_05588_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13584_ (.A1(_04400_),
    .A2(_05588_),
    .ZN(_05589_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13585_ (.A1(_05587_),
    .A2(_05589_),
    .Z(_05590_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13586_ (.A1(_05586_),
    .A2(_05590_),
    .ZN(_05591_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _13587_ (.A1(_04238_),
    .A2(_04945_),
    .B1(_05518_),
    .B2(_04847_),
    .ZN(_05592_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _13588_ (.A1(_04848_),
    .A2(_04850_),
    .A3(_04945_),
    .A4(_05518_),
    .ZN(_05593_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _13589_ (.A1(_05515_),
    .A2(_05592_),
    .B(_05593_),
    .ZN(_05594_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13590_ (.A1(_04476_),
    .A2(_05077_),
    .Z(_05595_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13591_ (.A1(_04236_),
    .A2(_04861_),
    .Z(_05596_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13592_ (.A1(_04220_),
    .A2(_04926_),
    .Z(_05597_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _13593_ (.A1(_05595_),
    .A2(_05596_),
    .A3(_05597_),
    .Z(_05598_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13594_ (.A1(_05594_),
    .A2(_05598_),
    .Z(_05599_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13595_ (.A1(_05591_),
    .A2(_05599_),
    .ZN(_05600_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13596_ (.A1(_05584_),
    .A2(_05600_),
    .ZN(_05601_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13597_ (.A1(_05582_),
    .A2(_05601_),
    .Z(_05602_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13598_ (.A1(_05477_),
    .A2(_05491_),
    .ZN(_05603_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _13599_ (.A1(net62),
    .A2(_05492_),
    .B(_05603_),
    .ZN(_05604_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13600_ (.A1(_05471_),
    .A2(_05472_),
    .Z(_05605_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _13601_ (.A1(_05471_),
    .A2(_05472_),
    .Z(_05606_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _13602_ (.A1(_05470_),
    .A2(_05605_),
    .B(_05606_),
    .ZN(_05607_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13603_ (.A1(_05479_),
    .A2(_05480_),
    .Z(_05608_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _13604_ (.A1(_05479_),
    .A2(_05480_),
    .Z(_05609_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13605_ (.A1(_05478_),
    .A2(_05608_),
    .B(_05609_),
    .ZN(_05610_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13606_ (.A1(_05158_),
    .A2(_05516_),
    .ZN(_05611_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13607_ (.A1(_04377_),
    .A2(_04751_),
    .ZN(_05612_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13608_ (.A1(_04317_),
    .A2(_04713_),
    .ZN(_05613_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _13609_ (.A1(_05611_),
    .A2(_05612_),
    .A3(_05613_),
    .Z(_05614_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13610_ (.A1(_05610_),
    .A2(_05614_),
    .ZN(_05615_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13611_ (.A1(_05607_),
    .A2(_05615_),
    .ZN(_05616_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13612_ (.A1(_05484_),
    .A2(_05489_),
    .ZN(_05617_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _13613_ (.A1(_05482_),
    .A2(_05490_),
    .B(_05617_),
    .ZN(_05618_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13614_ (.A1(_04864_),
    .A2(_04445_),
    .ZN(_05619_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _13615_ (.A1(_03364_),
    .A2(_04854_),
    .A3(_05220_),
    .ZN(_05620_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _13616_ (.A1(_03383_),
    .A2(_04342_),
    .A3(_04804_),
    .ZN(_05621_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13617_ (.A1(_05620_),
    .A2(_05621_),
    .Z(_05622_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13618_ (.A1(_05619_),
    .A2(_05622_),
    .Z(_05623_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _13619_ (.I(_05487_),
    .Z(_05624_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13620_ (.I(_05145_),
    .Z(_05625_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _13621_ (.I(_05625_),
    .Z(_05626_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _13622_ (.A1(_05231_),
    .A2(_05624_),
    .B1(_05626_),
    .B2(_04473_),
    .ZN(_05627_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _13623_ (.A1(_04473_),
    .A2(_05231_),
    .A3(_05624_),
    .A4(_05626_),
    .ZN(_05628_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _13624_ (.A1(_05485_),
    .A2(_05627_),
    .B(_05628_),
    .ZN(_05629_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _13625_ (.A1(_04485_),
    .A2(_04884_),
    .ZN(_05630_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _13626_ (.A1(_03316_),
    .A2(_04163_),
    .A3(_05208_),
    .ZN(_05631_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _13627_ (.A1(_03332_),
    .A2(_04522_),
    .A3(_05487_),
    .ZN(_05632_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _13628_ (.A1(_05630_),
    .A2(_05631_),
    .A3(_05632_),
    .ZN(_05633_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13629_ (.A1(_05629_),
    .A2(_05633_),
    .ZN(_05634_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13630_ (.A1(_05623_),
    .A2(_05634_),
    .Z(_05635_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13631_ (.A1(_05618_),
    .A2(_05635_),
    .ZN(_05636_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13632_ (.A1(_05616_),
    .A2(_05636_),
    .Z(_05637_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13633_ (.A1(_05604_),
    .A2(_05637_),
    .ZN(_05638_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13634_ (.A1(_05602_),
    .A2(_05638_),
    .Z(_05639_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13635_ (.A1(_05579_),
    .A2(_05639_),
    .Z(_05640_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13636_ (.A1(_05577_),
    .A2(_05640_),
    .Z(_05641_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _13637_ (.A1(_05555_),
    .A2(_05559_),
    .A3(_05641_),
    .ZN(_05642_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _13638_ (.A1(_05553_),
    .A2(_05642_),
    .ZN(_05643_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _13639_ (.A1(_05549_),
    .A2(_05550_),
    .A3(_05643_),
    .Z(_05644_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _13640_ (.A1(_05549_),
    .A2(_05550_),
    .B(_05643_),
    .ZN(_05645_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13641_ (.A1(_05644_),
    .A2(_05645_),
    .Z(_05646_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _13642_ (.I(\filters.low[1] ),
    .Z(_05647_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13643_ (.A1(_05647_),
    .A2(_03219_),
    .ZN(_05648_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _13644_ (.A1(_03251_),
    .A2(_03376_),
    .B(_05648_),
    .ZN(_05649_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13645_ (.A1(_05646_),
    .A2(_05649_),
    .Z(_05650_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13646_ (.A1(_05548_),
    .A2(_05650_),
    .Z(_05651_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13647_ (.A1(_05547_),
    .A2(_05651_),
    .ZN(_05652_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13648_ (.I(_01822_),
    .Z(_05653_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _13649_ (.A1(_03251_),
    .A2(_05545_),
    .B(_05652_),
    .C(_05653_),
    .ZN(_00527_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13650_ (.A1(_05527_),
    .A2(_05530_),
    .ZN(_05654_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13651_ (.A1(_05553_),
    .A2(_05642_),
    .ZN(_05655_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13652_ (.A1(_05553_),
    .A2(_05642_),
    .ZN(_05656_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _13653_ (.A1(_05654_),
    .A2(_05655_),
    .B(_05656_),
    .ZN(_05657_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _13654_ (.A1(net35),
    .A2(net40),
    .B(_05531_),
    .C(_05643_),
    .ZN(_05658_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _13655_ (.A1(_05568_),
    .A2(_05575_),
    .Z(_05659_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _13656_ (.A1(_05565_),
    .A2(_05576_),
    .B(_05659_),
    .ZN(_05660_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13657_ (.A1(_05579_),
    .A2(_05639_),
    .ZN(_05661_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _13658_ (.A1(_05577_),
    .A2(_05640_),
    .B(_05661_),
    .ZN(_05662_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13659_ (.I(_05570_),
    .Z(_05663_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13660_ (.A1(_04645_),
    .A2(_05663_),
    .A3(_05572_),
    .ZN(_05664_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13661_ (.A1(_04562_),
    .A2(_05561_),
    .A3(_05574_),
    .ZN(_05665_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13662_ (.A1(_05664_),
    .A2(_05665_),
    .Z(_05666_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13663_ (.A1(_05584_),
    .A2(_05600_),
    .ZN(_05667_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13664_ (.A1(_05582_),
    .A2(_05601_),
    .ZN(_05668_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13665_ (.A1(_05667_),
    .A2(_05668_),
    .ZN(_05669_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13666_ (.A1(_04500_),
    .A2(_05663_),
    .ZN(_05670_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13667_ (.I(_05585_),
    .Z(_05671_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13668_ (.A1(_04578_),
    .A2(_05671_),
    .A3(_05590_),
    .ZN(_05672_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13669_ (.A1(_05587_),
    .A2(_05589_),
    .B(_05672_),
    .ZN(_05673_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13670_ (.A1(_04211_),
    .A2(_05671_),
    .ZN(_05674_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13671_ (.A1(_05673_),
    .A2(_05674_),
    .ZN(_05675_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13672_ (.A1(_05670_),
    .A2(_05675_),
    .Z(_05676_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13673_ (.A1(_05669_),
    .A2(_05676_),
    .ZN(_05677_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13674_ (.A1(_05666_),
    .A2(_05677_),
    .Z(_05678_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13675_ (.I(_05602_),
    .ZN(_05679_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13676_ (.A1(_05604_),
    .A2(_05637_),
    .ZN(_05680_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13677_ (.A1(_05679_),
    .A2(_05638_),
    .B(_05680_),
    .ZN(_05681_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13678_ (.A1(_05594_),
    .A2(_05598_),
    .Z(_05682_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _13679_ (.A1(_05591_),
    .A2(_05599_),
    .B(_05682_),
    .ZN(_05683_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13680_ (.A1(_04512_),
    .A2(_04447_),
    .A3(_05481_),
    .ZN(_05684_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _13681_ (.A1(_05609_),
    .A2(_05684_),
    .B(_05614_),
    .ZN(_05685_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _13682_ (.A1(_05607_),
    .A2(_05615_),
    .B(_05685_),
    .ZN(_05686_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13683_ (.I(_05588_),
    .Z(_05687_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13684_ (.A1(_04176_),
    .A2(_05687_),
    .ZN(_05688_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13685_ (.A1(_04294_),
    .A2(_05260_),
    .ZN(_05689_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13686_ (.I0(\filters.high[22] ),
    .I1(\filters.band[22] ),
    .S(_05179_),
    .Z(_05690_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13687_ (.A1(_04400_),
    .A2(_05690_),
    .ZN(_05691_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13688_ (.A1(_05689_),
    .A2(_05691_),
    .Z(_05692_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13689_ (.A1(_05688_),
    .A2(_05692_),
    .ZN(_05693_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _13690_ (.A1(_05596_),
    .A2(_05597_),
    .Z(_05694_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13691_ (.A1(_05596_),
    .A2(_05597_),
    .Z(_05695_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _13692_ (.A1(_05595_),
    .A2(_05694_),
    .B(_05695_),
    .ZN(_05696_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13693_ (.A1(_04230_),
    .A2(_05256_),
    .ZN(_05697_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13694_ (.A1(_04694_),
    .A2(_05075_),
    .ZN(_05698_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13695_ (.A1(_04222_),
    .A2(_05280_),
    .ZN(_05699_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _13696_ (.A1(_05697_),
    .A2(_05698_),
    .A3(_05699_),
    .ZN(_05700_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _13697_ (.A1(_05693_),
    .A2(_05696_),
    .A3(_05700_),
    .Z(_05701_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13698_ (.A1(_05686_),
    .A2(_05701_),
    .ZN(_05702_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13699_ (.A1(_05683_),
    .A2(_05702_),
    .ZN(_05703_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13700_ (.A1(_05618_),
    .A2(_05635_),
    .ZN(_05704_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _13701_ (.A1(_05616_),
    .A2(_05636_),
    .B(_05704_),
    .ZN(_05705_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13702_ (.A1(_05612_),
    .A2(_05613_),
    .Z(_05706_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _13703_ (.A1(_05612_),
    .A2(_05613_),
    .Z(_05707_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _13704_ (.A1(_05611_),
    .A2(_05706_),
    .B(_05707_),
    .ZN(_05708_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13705_ (.A1(_05620_),
    .A2(_05621_),
    .Z(_05709_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _13706_ (.A1(_05620_),
    .A2(_05621_),
    .Z(_05710_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13707_ (.A1(_05619_),
    .A2(_05709_),
    .B(_05710_),
    .ZN(_05711_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13708_ (.A1(_04325_),
    .A2(_04924_),
    .ZN(_05712_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13709_ (.A1(_04452_),
    .A2(_04713_),
    .ZN(_05713_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13710_ (.A1(_04449_),
    .A2(_04945_),
    .ZN(_05714_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _13711_ (.A1(_05712_),
    .A2(_05713_),
    .A3(_05714_),
    .Z(_05715_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13712_ (.A1(_05711_),
    .A2(_05715_),
    .ZN(_05716_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13713_ (.A1(_05708_),
    .A2(_05716_),
    .ZN(_05717_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13714_ (.A1(_05629_),
    .A2(_05633_),
    .ZN(_05718_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13715_ (.A1(_05623_),
    .A2(_05634_),
    .B(_05718_),
    .ZN(_05719_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13716_ (.A1(_04802_),
    .A2(_04753_),
    .ZN(_05720_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _13717_ (.I(_04825_),
    .Z(_05721_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _13718_ (.A1(_03383_),
    .A2(_04342_),
    .A3(_05721_),
    .ZN(_05722_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _13719_ (.A1(_03398_),
    .A2(_04403_),
    .A3(_04805_),
    .ZN(_05723_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13720_ (.A1(_05722_),
    .A2(_05723_),
    .Z(_05724_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13721_ (.A1(_05720_),
    .A2(_05724_),
    .Z(_05725_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13722_ (.A1(_05631_),
    .A2(_05632_),
    .Z(_05726_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _13723_ (.A1(_05631_),
    .A2(_05632_),
    .Z(_05727_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _13724_ (.A1(_05630_),
    .A2(_05726_),
    .B(_05727_),
    .ZN(_05728_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13725_ (.A1(_04274_),
    .A2(_04819_),
    .Z(_05729_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _13726_ (.A1(_03333_),
    .A2(_04522_),
    .A3(_05625_),
    .ZN(_05730_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _13727_ (.I(_04881_),
    .Z(_05731_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _13728_ (.I(_05731_),
    .Z(_05732_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13729_ (.A1(_03350_),
    .A2(_04192_),
    .A3(_05732_),
    .ZN(_05733_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13730_ (.A1(_05730_),
    .A2(_05733_),
    .Z(_05734_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13731_ (.A1(_05729_),
    .A2(_05734_),
    .Z(_05735_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13732_ (.A1(_05728_),
    .A2(_05735_),
    .ZN(_05736_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13733_ (.A1(_05725_),
    .A2(_05736_),
    .Z(_05737_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13734_ (.A1(_05719_),
    .A2(_05737_),
    .ZN(_05738_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13735_ (.A1(_05717_),
    .A2(_05738_),
    .Z(_05739_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _13736_ (.A1(_05703_),
    .A2(_05705_),
    .A3(_05739_),
    .ZN(_05740_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _13737_ (.A1(_05678_),
    .A2(_05681_),
    .A3(_05740_),
    .ZN(_05741_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _13738_ (.A1(_05662_),
    .A2(_05741_),
    .Z(_05742_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _13739_ (.A1(_05660_),
    .A2(_05742_),
    .Z(_05743_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13740_ (.A1(_05559_),
    .A2(_05641_),
    .ZN(_05744_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13741_ (.A1(_05559_),
    .A2(_05641_),
    .ZN(_05745_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _13742_ (.A1(_05555_),
    .A2(_05744_),
    .B(_05745_),
    .ZN(_05746_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _13743_ (.A1(_05743_),
    .A2(_05746_),
    .Z(_05747_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13744_ (.A1(_05657_),
    .A2(_05658_),
    .B(_05747_),
    .ZN(_05748_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _13745_ (.A1(_05747_),
    .A2(_05657_),
    .A3(_05658_),
    .Z(_05749_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13746_ (.A1(_05748_),
    .A2(_05749_),
    .ZN(_05750_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _13747_ (.I(_05750_),
    .Z(_05751_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _13748_ (.I(_05751_),
    .Z(_05752_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13749_ (.A1(_03268_),
    .A2(_03375_),
    .ZN(_05753_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13750_ (.A1(_03269_),
    .A2(_03346_),
    .B(_05753_),
    .ZN(_05754_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13751_ (.I(_05754_),
    .Z(_05755_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _13752_ (.A1(_05644_),
    .A2(_05645_),
    .B(_05649_),
    .ZN(_05756_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13753_ (.A1(_05644_),
    .A2(_05645_),
    .A3(_05649_),
    .ZN(_05757_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _13754_ (.A1(_05537_),
    .A2(_05756_),
    .B(_05757_),
    .ZN(_05758_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _13755_ (.A1(_05752_),
    .A2(_05755_),
    .A3(_05758_),
    .Z(_05759_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13756_ (.A1(_05547_),
    .A2(_05759_),
    .ZN(_05760_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _13757_ (.A1(_03269_),
    .A2(_05545_),
    .B(_05760_),
    .C(_05653_),
    .ZN(_00528_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _13758_ (.A1(_05669_),
    .A2(_05676_),
    .Z(_05761_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _13759_ (.A1(_05666_),
    .A2(_05677_),
    .B(_05761_),
    .ZN(_05762_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _13760_ (.A1(_05681_),
    .A2(_05740_),
    .Z(_05763_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13761_ (.A1(_05681_),
    .A2(_05740_),
    .Z(_05764_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _13762_ (.A1(_05678_),
    .A2(_05763_),
    .B(_05764_),
    .ZN(_05765_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13763_ (.I(_05671_),
    .Z(_05766_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13764_ (.A1(_04667_),
    .A2(_05766_),
    .A3(_05673_),
    .ZN(_05767_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13765_ (.A1(_05563_),
    .A2(_05663_),
    .A3(_05675_),
    .ZN(_05768_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13766_ (.A1(_05767_),
    .A2(_05768_),
    .Z(_05769_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13767_ (.A1(_05686_),
    .A2(_05701_),
    .ZN(_05770_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13768_ (.A1(_05683_),
    .A2(_05702_),
    .ZN(_05771_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13769_ (.A1(_05770_),
    .A2(_05771_),
    .ZN(_05772_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13770_ (.A1(_04630_),
    .A2(_05766_),
    .ZN(_05773_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13771_ (.I(_05687_),
    .Z(_05774_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13772_ (.I(_05774_),
    .Z(_05775_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13773_ (.A1(_04597_),
    .A2(_05775_),
    .A3(_05692_),
    .ZN(_05776_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13774_ (.A1(_05689_),
    .A2(_05691_),
    .B(_05776_),
    .ZN(_05777_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13775_ (.A1(_04764_),
    .A2(_05775_),
    .ZN(_05778_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13776_ (.A1(_05777_),
    .A2(_05778_),
    .ZN(_05779_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13777_ (.A1(_05773_),
    .A2(_05779_),
    .Z(_05780_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13778_ (.A1(_05772_),
    .A2(_05780_),
    .ZN(_05781_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13779_ (.A1(_05769_),
    .A2(_05781_),
    .Z(_05782_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13780_ (.A1(_05705_),
    .A2(_05739_),
    .ZN(_05783_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13781_ (.A1(_05705_),
    .A2(_05739_),
    .ZN(_05784_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13782_ (.A1(_05703_),
    .A2(_05783_),
    .B(_05784_),
    .ZN(_05785_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13783_ (.I(_05700_),
    .ZN(_05786_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13784_ (.A1(_05696_),
    .A2(_05786_),
    .ZN(_05787_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13785_ (.A1(_05696_),
    .A2(_05786_),
    .ZN(_05788_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _13786_ (.A1(_05693_),
    .A2(_05787_),
    .B(_05788_),
    .ZN(_05789_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13787_ (.A1(_04966_),
    .A2(_04447_),
    .A3(_05622_),
    .ZN(_05790_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _13788_ (.A1(_05710_),
    .A2(_05790_),
    .B(_05715_),
    .ZN(_05791_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _13789_ (.A1(_05708_),
    .A2(_05716_),
    .B(_05791_),
    .ZN(_05792_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13790_ (.I(_05690_),
    .Z(_05793_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13791_ (.A1(_04525_),
    .A2(_05793_),
    .ZN(_05794_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13792_ (.A1(_04200_),
    .A2(_05500_),
    .ZN(_05795_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13793_ (.I0(\filters.high[23] ),
    .I1(\filters.band[23] ),
    .S(_03187_),
    .Z(_05796_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13794_ (.A1(_04487_),
    .A2(_05796_),
    .ZN(_05797_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13795_ (.A1(_05795_),
    .A2(_05797_),
    .Z(_05798_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13796_ (.A1(_05794_),
    .A2(_05798_),
    .ZN(_05799_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13797_ (.I(_04471_),
    .Z(_05800_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _13798_ (.A1(_05512_),
    .A2(_05091_),
    .B1(_05079_),
    .B2(_05800_),
    .ZN(_05801_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _13799_ (.A1(_04694_),
    .A2(_05800_),
    .A3(_05091_),
    .A4(_05079_),
    .ZN(_05802_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _13800_ (.A1(_05697_),
    .A2(_05801_),
    .B(_05802_),
    .ZN(_05803_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13801_ (.A1(_04705_),
    .A2(_05260_),
    .ZN(_05804_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13802_ (.A1(_04728_),
    .A2(_05078_),
    .ZN(_05805_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13803_ (.A1(_04221_),
    .A2(_05187_),
    .ZN(_05806_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _13804_ (.A1(_05804_),
    .A2(_05805_),
    .A3(_05806_),
    .ZN(_05807_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13805_ (.A1(_05803_),
    .A2(_05807_),
    .Z(_05808_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13806_ (.A1(_05799_),
    .A2(_05808_),
    .ZN(_05809_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13807_ (.A1(_05792_),
    .A2(_05809_),
    .ZN(_05810_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13808_ (.A1(_05789_),
    .A2(_05810_),
    .Z(_05811_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13809_ (.A1(_05719_),
    .A2(_05737_),
    .ZN(_05812_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _13810_ (.A1(_05717_),
    .A2(_05738_),
    .B(_05812_),
    .ZN(_05813_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13811_ (.A1(_05713_),
    .A2(_05714_),
    .Z(_05814_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _13812_ (.A1(_05713_),
    .A2(_05714_),
    .Z(_05815_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _13813_ (.A1(_05712_),
    .A2(_05814_),
    .B(_05815_),
    .ZN(_05816_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13814_ (.A1(_05722_),
    .A2(_05723_),
    .Z(_05817_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _13815_ (.A1(_05722_),
    .A2(_05723_),
    .Z(_05818_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13816_ (.A1(_05720_),
    .A2(_05817_),
    .B(_05818_),
    .ZN(_05819_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13817_ (.A1(_05158_),
    .A2(_05074_),
    .Z(_05820_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13818_ (.A1(_04451_),
    .A2(_05516_),
    .ZN(_05821_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13819_ (.A1(_04893_),
    .A2(_05518_),
    .ZN(_05822_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _13820_ (.A1(_05820_),
    .A2(_05821_),
    .A3(_05822_),
    .ZN(_05823_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13821_ (.A1(_05819_),
    .A2(_05823_),
    .ZN(_05824_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13822_ (.A1(_05816_),
    .A2(_05824_),
    .ZN(_05825_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13823_ (.A1(_05728_),
    .A2(_05735_),
    .ZN(_05826_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13824_ (.A1(_05725_),
    .A2(_05736_),
    .B(_05826_),
    .ZN(_05827_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13825_ (.I(_05469_),
    .Z(_05828_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13826_ (.A1(_04445_),
    .A2(_05828_),
    .ZN(_05829_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13827_ (.A1(_04864_),
    .A2(_05721_),
    .ZN(_05830_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13828_ (.A1(_04753_),
    .A2(_05466_),
    .ZN(_05831_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _13829_ (.A1(_05829_),
    .A2(_05830_),
    .A3(_05831_),
    .Z(_05832_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13830_ (.A1(_05730_),
    .A2(_05733_),
    .ZN(_05833_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _13831_ (.A1(_05729_),
    .A2(_05734_),
    .B(_05833_),
    .ZN(_05834_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13832_ (.A1(_04397_),
    .A2(_04818_),
    .Z(_05835_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _13833_ (.A1(_03349_),
    .A2(_04191_),
    .A3(_05145_),
    .ZN(_05836_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13834_ (.A1(_03363_),
    .A2(_04854_),
    .A3(_05731_),
    .ZN(_05837_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13835_ (.A1(_05836_),
    .A2(_05837_),
    .Z(_05838_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13836_ (.A1(_05835_),
    .A2(_05838_),
    .ZN(_05839_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13837_ (.A1(_05834_),
    .A2(_05839_),
    .ZN(_05840_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13838_ (.A1(_05832_),
    .A2(_05840_),
    .Z(_05841_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13839_ (.A1(_05827_),
    .A2(_05841_),
    .ZN(_05842_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13840_ (.A1(_05825_),
    .A2(_05842_),
    .Z(_05843_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _13841_ (.A1(_05811_),
    .A2(_05813_),
    .A3(_05843_),
    .Z(_05844_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _13842_ (.A1(_05782_),
    .A2(_05785_),
    .A3(_05844_),
    .ZN(_05845_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _13843_ (.A1(_05762_),
    .A2(_05765_),
    .A3(_05845_),
    .ZN(_05846_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13844_ (.A1(_05662_),
    .A2(_05741_),
    .ZN(_05847_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _13845_ (.A1(_05660_),
    .A2(_05742_),
    .B(_05847_),
    .ZN(_05848_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _13846_ (.A1(_05846_),
    .A2(_05848_),
    .Z(_05849_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13847_ (.A1(_05743_),
    .A2(_05746_),
    .ZN(_05850_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13848_ (.A1(_05850_),
    .A2(_05748_),
    .ZN(_05851_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _13849_ (.A1(_05849_),
    .A2(_05851_),
    .ZN(_05852_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13850_ (.I(_03376_),
    .Z(_05853_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13851_ (.A1(_03282_),
    .A2(_03220_),
    .ZN(_05854_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _13852_ (.A1(_03284_),
    .A2(_05853_),
    .B(_05854_),
    .ZN(_05855_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13853_ (.A1(_05852_),
    .A2(_05855_),
    .Z(_05856_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13854_ (.A1(_05752_),
    .A2(_05755_),
    .ZN(_05857_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13855_ (.A1(_05548_),
    .A2(_05650_),
    .ZN(_05858_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13856_ (.A1(_05757_),
    .A2(_05858_),
    .Z(_05859_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13857_ (.A1(_05752_),
    .A2(_05755_),
    .ZN(_05860_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13858_ (.A1(_05857_),
    .A2(_05859_),
    .B(_05860_),
    .ZN(_05861_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13859_ (.A1(_05856_),
    .A2(_05861_),
    .Z(_05862_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13860_ (.A1(_05547_),
    .A2(_05862_),
    .ZN(_05863_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _13861_ (.A1(_03284_),
    .A2(_05545_),
    .B(_05863_),
    .C(_05653_),
    .ZN(_00529_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _13862_ (.A1(_05852_),
    .A2(_05855_),
    .ZN(_05864_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _13863_ (.A1(_05750_),
    .A2(_05755_),
    .Z(_05865_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13864_ (.A1(_05750_),
    .A2(_05754_),
    .Z(_05866_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _13865_ (.A1(_05865_),
    .A2(_05758_),
    .B(_05866_),
    .ZN(_05867_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13866_ (.A1(_05852_),
    .A2(_05855_),
    .ZN(_05868_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _13867_ (.A1(_05864_),
    .A2(_05867_),
    .B(_05868_),
    .ZN(_05869_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13868_ (.A1(_05531_),
    .A2(_05643_),
    .ZN(_05870_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _13869_ (.A1(_05747_),
    .A2(_05870_),
    .A3(_05849_),
    .ZN(_05871_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _13870_ (.A1(_05747_),
    .A2(_05657_),
    .A3(_05849_),
    .ZN(_05872_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13871_ (.A1(_05743_),
    .A2(_05746_),
    .Z(_05873_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13872_ (.A1(_05846_),
    .A2(_05848_),
    .ZN(_05874_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13873_ (.A1(_05846_),
    .A2(_05848_),
    .ZN(_05875_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _13874_ (.A1(_05873_),
    .A2(_05874_),
    .B(_05875_),
    .ZN(_05876_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _13875_ (.A1(_05432_),
    .A2(_05871_),
    .B(_05872_),
    .C(_05876_),
    .ZN(_05877_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _13876_ (.A1(_05772_),
    .A2(_05780_),
    .Z(_05878_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _13877_ (.A1(_05769_),
    .A2(_05781_),
    .B(_05878_),
    .ZN(_05879_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _13878_ (.A1(_05785_),
    .A2(_05844_),
    .Z(_05880_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13879_ (.A1(_05785_),
    .A2(_05844_),
    .Z(_05881_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _13880_ (.A1(_05782_),
    .A2(_05880_),
    .B(_05881_),
    .ZN(_05882_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13881_ (.I(_05775_),
    .Z(_05883_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13882_ (.A1(_04667_),
    .A2(_05883_),
    .A3(_05777_),
    .ZN(_05884_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13883_ (.A1(_05440_),
    .A2(_05766_),
    .A3(_05779_),
    .ZN(_05885_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13884_ (.A1(_05884_),
    .A2(_05885_),
    .Z(_05886_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13885_ (.A1(_05792_),
    .A2(_05809_),
    .ZN(_05887_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13886_ (.A1(_05789_),
    .A2(_05810_),
    .ZN(_05888_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13887_ (.A1(_05887_),
    .A2(_05888_),
    .ZN(_05889_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13888_ (.A1(_04561_),
    .A2(_05883_),
    .ZN(_05890_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13889_ (.I(_05793_),
    .Z(_05891_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13890_ (.I(_05891_),
    .Z(_05892_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13891_ (.A1(_04597_),
    .A2(_05892_),
    .A3(_05798_),
    .ZN(_05893_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13892_ (.A1(_05795_),
    .A2(_05797_),
    .B(_05893_),
    .ZN(_05894_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13893_ (.A1(_04642_),
    .A2(_05892_),
    .ZN(_05895_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13894_ (.A1(_05894_),
    .A2(_05895_),
    .ZN(_05896_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13895_ (.A1(_05890_),
    .A2(_05896_),
    .Z(_05897_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13896_ (.A1(_05889_),
    .A2(_05897_),
    .ZN(_05898_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13897_ (.A1(_05886_),
    .A2(_05898_),
    .Z(_05899_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13898_ (.I(_05811_),
    .ZN(_05900_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13899_ (.A1(_05813_),
    .A2(_05843_),
    .ZN(_05901_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13900_ (.A1(_05813_),
    .A2(_05843_),
    .ZN(_05902_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13901_ (.A1(_05900_),
    .A2(_05901_),
    .B(_05902_),
    .ZN(_05903_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13902_ (.A1(_05827_),
    .A2(_05841_),
    .ZN(_05904_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _13903_ (.A1(_05825_),
    .A2(_05842_),
    .B(_05904_),
    .ZN(_05905_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13904_ (.A1(_05821_),
    .A2(_05822_),
    .ZN(_05906_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13905_ (.A1(_05821_),
    .A2(_05822_),
    .ZN(_05907_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _13906_ (.A1(_05820_),
    .A2(_05906_),
    .B(_05907_),
    .ZN(_05908_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13907_ (.I(_05229_),
    .Z(_05909_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _13908_ (.A1(_04406_),
    .A2(_05909_),
    .B1(_05466_),
    .B2(_04929_),
    .ZN(_05910_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _13909_ (.A1(_04406_),
    .A2(_04929_),
    .A3(_05465_),
    .A4(_05466_),
    .ZN(_05911_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _13910_ (.A1(_05829_),
    .A2(_05910_),
    .B(_05911_),
    .ZN(_05912_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13911_ (.A1(_04324_),
    .A2(_05078_),
    .Z(_05913_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13912_ (.A1(_04451_),
    .A2(_04862_),
    .ZN(_05914_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13913_ (.A1(_04317_),
    .A2(_04927_),
    .ZN(_05915_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _13914_ (.A1(_05913_),
    .A2(_05914_),
    .A3(_05915_),
    .Z(_05916_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13915_ (.A1(_05912_),
    .A2(_05916_),
    .ZN(_05917_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13916_ (.A1(_05908_),
    .A2(_05917_),
    .ZN(_05918_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _13917_ (.A1(_05834_),
    .A2(_05839_),
    .Z(_05919_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _13918_ (.A1(_05832_),
    .A2(_05840_),
    .B(_05919_),
    .ZN(_05920_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13919_ (.A1(_05836_),
    .A2(_05837_),
    .ZN(_05921_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _13920_ (.A1(_05835_),
    .A2(_05838_),
    .B(_05921_),
    .ZN(_05922_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13921_ (.A1(_04272_),
    .A2(_05208_),
    .ZN(_05923_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13922_ (.A1(_04396_),
    .A2(_05731_),
    .ZN(_05924_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13923_ (.A1(_04483_),
    .A2(_04818_),
    .ZN(_05925_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _13924_ (.A1(_05923_),
    .A2(_05924_),
    .A3(_05925_),
    .Z(_05926_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13925_ (.A1(_05922_),
    .A2(_05926_),
    .ZN(_05927_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13926_ (.A1(_04801_),
    .A2(_05183_),
    .ZN(_05928_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13927_ (.A1(_04752_),
    .A2(_05229_),
    .ZN(_05929_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _13928_ (.I(_05230_),
    .Z(_05930_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13929_ (.A1(_05828_),
    .A2(_05930_),
    .ZN(_05931_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _13930_ (.A1(_05928_),
    .A2(_05929_),
    .A3(_05931_),
    .Z(_05932_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13931_ (.A1(_05927_),
    .A2(_05932_),
    .Z(_05933_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13932_ (.A1(_05920_),
    .A2(_05933_),
    .ZN(_05934_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _13933_ (.A1(_05918_),
    .A2(_05934_),
    .Z(_05935_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13934_ (.A1(_05803_),
    .A2(_05807_),
    .Z(_05936_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _13935_ (.A1(_05799_),
    .A2(_05808_),
    .B(_05936_),
    .ZN(_05937_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13936_ (.A1(_04446_),
    .A2(_04766_),
    .A3(_05724_),
    .ZN(_05938_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _13937_ (.A1(_05818_),
    .A2(_05938_),
    .B(_05823_),
    .ZN(_05939_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _13938_ (.A1(_05816_),
    .A2(_05824_),
    .B(_05939_),
    .ZN(_05940_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13939_ (.A1(_04176_),
    .A2(_05796_),
    .ZN(_05941_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13940_ (.A1(_04294_),
    .A2(_05504_),
    .ZN(_05942_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13941_ (.I0(\filters.high[24] ),
    .I1(\filters.band[24] ),
    .S(_05179_),
    .Z(_05943_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13942_ (.A1(_04186_),
    .A2(_05943_),
    .ZN(_05944_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13943_ (.A1(_05942_),
    .A2(_05944_),
    .Z(_05945_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13944_ (.A1(_05941_),
    .A2(_05945_),
    .ZN(_05946_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _13945_ (.I(_05186_),
    .Z(_05947_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _13946_ (.A1(_04238_),
    .A2(_05279_),
    .B1(_05947_),
    .B2(_04847_),
    .ZN(_05948_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _13947_ (.A1(_04238_),
    .A2(_04847_),
    .A3(_05279_),
    .A4(_05947_),
    .ZN(_05949_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _13948_ (.A1(_05804_),
    .A2(_05948_),
    .B(_05949_),
    .ZN(_05950_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13949_ (.A1(_04229_),
    .A2(_05351_),
    .ZN(_05951_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13950_ (.A1(_04254_),
    .A2(_05185_),
    .ZN(_05952_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13951_ (.A1(_04392_),
    .A2(_05347_),
    .ZN(_05953_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _13952_ (.A1(_05951_),
    .A2(_05952_),
    .A3(_05953_),
    .ZN(_05954_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13953_ (.A1(_05950_),
    .A2(_05954_),
    .Z(_05955_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13954_ (.A1(_05946_),
    .A2(_05955_),
    .ZN(_05956_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13955_ (.A1(_05940_),
    .A2(_05956_),
    .ZN(_05957_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13956_ (.A1(_05937_),
    .A2(_05957_),
    .ZN(_05958_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _13957_ (.A1(_05905_),
    .A2(_05935_),
    .A3(_05958_),
    .ZN(_05959_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _13958_ (.A1(_05903_),
    .A2(_05959_),
    .Z(_05960_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13959_ (.A1(_05899_),
    .A2(_05960_),
    .ZN(_05961_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _13960_ (.A1(_05882_),
    .A2(_05961_),
    .Z(_05962_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13961_ (.A1(_05879_),
    .A2(_05962_),
    .ZN(_05963_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13962_ (.A1(_05765_),
    .A2(_05845_),
    .ZN(_05964_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13963_ (.A1(_05765_),
    .A2(_05845_),
    .ZN(_05965_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _13964_ (.A1(_05762_),
    .A2(_05964_),
    .B(_05965_),
    .ZN(_05966_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _13965_ (.A1(_05966_),
    .A2(_05963_),
    .Z(_05967_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _13966_ (.A1(_05877_),
    .A2(_05967_),
    .Z(_05968_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _13967_ (.I(\filters.low[4] ),
    .Z(_05969_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _13968_ (.A1(_05969_),
    .A2(_03471_),
    .ZN(_05970_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _13969_ (.A1(_03299_),
    .A2(_03471_),
    .B(_05970_),
    .ZN(_05971_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13970_ (.A1(_05968_),
    .A2(_05971_),
    .Z(_05972_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13971_ (.A1(_05869_),
    .A2(_05972_),
    .Z(_05973_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13972_ (.A1(\filters.band[4] ),
    .A2(_05540_),
    .B(_05541_),
    .ZN(_05974_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _13973_ (.A1(_04161_),
    .A2(_05973_),
    .B(_05974_),
    .ZN(_00530_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13974_ (.I(_05543_),
    .Z(_05975_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _13975_ (.A1(_05889_),
    .A2(_05897_),
    .Z(_05976_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _13976_ (.A1(_05886_),
    .A2(_05898_),
    .B(_05976_),
    .ZN(_05977_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13977_ (.A1(_05903_),
    .A2(_05959_),
    .Z(_05978_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _13978_ (.A1(_05899_),
    .A2(_05960_),
    .B(_05978_),
    .ZN(_05979_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13979_ (.I(_05892_),
    .Z(_05980_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13980_ (.A1(_05560_),
    .A2(_05980_),
    .A3(_05894_),
    .ZN(_05981_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _13981_ (.I(_04631_),
    .Z(_05982_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13982_ (.A1(_05982_),
    .A2(_05883_),
    .A3(_05896_),
    .ZN(_05983_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13983_ (.A1(_05981_),
    .A2(_05983_),
    .Z(_05984_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13984_ (.A1(_05940_),
    .A2(_05956_),
    .ZN(_05985_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13985_ (.A1(_05937_),
    .A2(_05957_),
    .ZN(_05986_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13986_ (.A1(_05985_),
    .A2(_05986_),
    .ZN(_05987_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13987_ (.A1(_04630_),
    .A2(_05892_),
    .ZN(_05988_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13988_ (.I(_05796_),
    .Z(_05989_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13989_ (.I(_05989_),
    .Z(_05990_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13990_ (.A1(_04616_),
    .A2(_05990_),
    .A3(_05945_),
    .ZN(_05991_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13991_ (.A1(_05942_),
    .A2(_05944_),
    .B(_05991_),
    .ZN(_05992_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13992_ (.A1(_04498_),
    .A2(_05990_),
    .ZN(_05993_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13993_ (.A1(_05992_),
    .A2(_05993_),
    .ZN(_05994_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13994_ (.A1(_05988_),
    .A2(_05994_),
    .Z(_05995_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13995_ (.A1(_05987_),
    .A2(_05995_),
    .ZN(_05996_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13996_ (.A1(_05984_),
    .A2(_05996_),
    .Z(_05997_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13997_ (.A1(_05905_),
    .A2(_05935_),
    .ZN(_05998_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13998_ (.A1(_05905_),
    .A2(_05935_),
    .ZN(_05999_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13999_ (.A1(_05998_),
    .A2(_05958_),
    .B(_05999_),
    .ZN(_06000_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _14000_ (.A1(_05950_),
    .A2(_05954_),
    .Z(_06001_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _14001_ (.A1(_05946_),
    .A2(_05955_),
    .B(_06001_),
    .ZN(_06002_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14002_ (.A1(_05912_),
    .A2(_05916_),
    .ZN(_06003_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _14003_ (.A1(_05908_),
    .A2(_05917_),
    .B(_06003_),
    .ZN(_06004_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _14004_ (.I(_05943_),
    .Z(_06005_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14005_ (.A1(_04529_),
    .A2(_06005_),
    .ZN(_06006_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14006_ (.A1(_04742_),
    .A2(_05588_),
    .ZN(_06007_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _14007_ (.I0(\filters.high[25] ),
    .I1(\filters.band[25] ),
    .S(_03187_),
    .Z(_06008_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14008_ (.A1(_04487_),
    .A2(_06008_),
    .ZN(_06009_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14009_ (.A1(_06007_),
    .A2(_06009_),
    .Z(_06010_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _14010_ (.A1(_06006_),
    .A2(_06010_),
    .ZN(_06011_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _14011_ (.A1(_05512_),
    .A2(_05256_),
    .B1(_05448_),
    .B2(_05800_),
    .ZN(_06012_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _14012_ (.A1(_04694_),
    .A2(_05800_),
    .A3(_05256_),
    .A4(_05447_),
    .ZN(_06013_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _14013_ (.A1(_05951_),
    .A2(_06012_),
    .B(_06013_),
    .ZN(_06014_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14014_ (.A1(_04728_),
    .A2(_05347_),
    .ZN(_06015_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14015_ (.A1(_04259_),
    .A2(_05351_),
    .ZN(_06016_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14016_ (.A1(_04230_),
    .A2(_05505_),
    .ZN(_06017_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _14017_ (.A1(_06015_),
    .A2(_06016_),
    .A3(_06017_),
    .ZN(_06018_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14018_ (.A1(_06014_),
    .A2(_06018_),
    .Z(_06019_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14019_ (.A1(_06011_),
    .A2(_06019_),
    .Z(_06020_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _14020_ (.A1(_06004_),
    .A2(_06020_),
    .ZN(_06021_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _14021_ (.A1(_06002_),
    .A2(_06021_),
    .ZN(_06022_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14022_ (.A1(_05920_),
    .A2(_05933_),
    .ZN(_06023_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _14023_ (.A1(_05918_),
    .A2(_05934_),
    .B(_06023_),
    .ZN(_06024_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _14024_ (.A1(_05922_),
    .A2(_05926_),
    .Z(_06025_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _14025_ (.A1(_05927_),
    .A2(_05932_),
    .B(_06025_),
    .ZN(_06026_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _14026_ (.I(_05625_),
    .Z(_06027_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _14027_ (.A1(_04397_),
    .A2(_05732_),
    .B1(_06027_),
    .B2(_04290_),
    .ZN(_06028_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _14028_ (.A1(_04290_),
    .A2(_04397_),
    .A3(_05732_),
    .A4(_06027_),
    .ZN(_06029_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _14029_ (.A1(_06028_),
    .A2(_05925_),
    .B(_06029_),
    .ZN(_06030_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14030_ (.A1(_03382_),
    .A2(_04341_),
    .A3(_05107_),
    .ZN(_06031_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14031_ (.A1(_03397_),
    .A2(_04403_),
    .A3(_04881_),
    .ZN(_06032_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _14032_ (.A1(_06031_),
    .A2(_06032_),
    .ZN(_06033_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14033_ (.A1(_04750_),
    .A2(_04884_),
    .ZN(_06034_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14034_ (.A1(_06033_),
    .A2(_06034_),
    .Z(_06035_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _14035_ (.A1(_06030_),
    .A2(_06035_),
    .ZN(_06036_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14036_ (.A1(_04801_),
    .A2(_04923_),
    .ZN(_06037_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14037_ (.A1(_05469_),
    .A2(_04825_),
    .ZN(_06038_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14038_ (.A1(_05516_),
    .A2(_05230_),
    .ZN(_06039_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _14039_ (.A1(_06037_),
    .A2(_06038_),
    .A3(_06039_),
    .Z(_06040_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14040_ (.A1(_06036_),
    .A2(_06040_),
    .Z(_06041_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _14041_ (.A1(_06026_),
    .A2(_06041_),
    .Z(_06042_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14042_ (.A1(_05914_),
    .A2(_05915_),
    .ZN(_06043_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14043_ (.A1(_05914_),
    .A2(_05915_),
    .ZN(_06044_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _14044_ (.A1(_05913_),
    .A2(_06043_),
    .B(_06044_),
    .ZN(_06045_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _14045_ (.A1(_04929_),
    .A2(_05465_),
    .B1(_05930_),
    .B2(_05828_),
    .ZN(_06046_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _14046_ (.A1(_04752_),
    .A2(_05828_),
    .A3(_05721_),
    .A4(_05930_),
    .ZN(_06047_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _14047_ (.A1(_05928_),
    .A2(_06046_),
    .B(_06047_),
    .ZN(_06048_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14048_ (.A1(_04377_),
    .A2(_05074_),
    .ZN(_06049_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14049_ (.A1(_04372_),
    .A2(_05078_),
    .ZN(_06050_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14050_ (.A1(_04325_),
    .A2(_05947_),
    .ZN(_06051_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _14051_ (.A1(_06049_),
    .A2(_06050_),
    .A3(_06051_),
    .Z(_06052_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14052_ (.A1(_06048_),
    .A2(_06052_),
    .Z(_06053_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14053_ (.A1(_06045_),
    .A2(_06053_),
    .Z(_06054_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _14054_ (.A1(_06042_),
    .A2(_06054_),
    .Z(_06055_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _14055_ (.A1(_06024_),
    .A2(_06055_),
    .ZN(_06056_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14056_ (.A1(_06022_),
    .A2(_06056_),
    .Z(_06057_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _14057_ (.A1(_05997_),
    .A2(_06000_),
    .A3(_06057_),
    .ZN(_06058_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _14058_ (.A1(_05977_),
    .A2(_05979_),
    .A3(_06058_),
    .ZN(_06059_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14059_ (.A1(_05882_),
    .A2(_05961_),
    .ZN(_06060_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _14060_ (.A1(_05879_),
    .A2(_05962_),
    .B(_06060_),
    .ZN(_06061_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _14061_ (.A1(_06059_),
    .A2(_06061_),
    .Z(_06062_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _14062_ (.A1(_05966_),
    .A2(_05963_),
    .ZN(_06063_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _14063_ (.A1(_05877_),
    .A2(_05967_),
    .B(net46),
    .ZN(_06064_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _14064_ (.A1(_06062_),
    .A2(_06064_),
    .Z(_06065_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _14065_ (.I(_03375_),
    .Z(_06066_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _14066_ (.I(_06066_),
    .Z(_06067_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14067_ (.A1(_03310_),
    .A2(_03377_),
    .ZN(_06068_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _14068_ (.A1(_03314_),
    .A2(_06067_),
    .B(_06068_),
    .ZN(_06069_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _14069_ (.A1(_06065_),
    .A2(_06069_),
    .ZN(_06070_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _14070_ (.A1(_06065_),
    .A2(_06069_),
    .Z(_06071_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14071_ (.A1(_06070_),
    .A2(_06071_),
    .ZN(_06072_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _14072_ (.I(_03472_),
    .Z(_06073_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _14073_ (.A1(_03299_),
    .A2(_06073_),
    .B(_05968_),
    .C(_05970_),
    .ZN(_06074_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14074_ (.A1(_05856_),
    .A2(_05861_),
    .ZN(_06075_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _14075_ (.A1(_05868_),
    .A2(_06075_),
    .B(_05972_),
    .ZN(_06076_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14076_ (.A1(_06074_),
    .A2(_06076_),
    .ZN(_06077_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _14077_ (.A1(_06072_),
    .A2(_06077_),
    .ZN(_06078_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14078_ (.A1(_05975_),
    .A2(_06078_),
    .ZN(_06079_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _14079_ (.A1(_03314_),
    .A2(_05545_),
    .B(_06079_),
    .C(_05653_),
    .ZN(_00531_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _14080_ (.I(_05544_),
    .Z(_06080_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _14081_ (.A1(_05987_),
    .A2(_05995_),
    .Z(_06081_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _14082_ (.A1(_05984_),
    .A2(_05996_),
    .B(_06081_),
    .ZN(_06082_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _14083_ (.A1(_06000_),
    .A2(_06057_),
    .Z(_06083_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _14084_ (.A1(_06000_),
    .A2(_06057_),
    .Z(_06084_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _14085_ (.A1(_05997_),
    .A2(_06083_),
    .B(_06084_),
    .ZN(_06085_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14086_ (.I(_05990_),
    .Z(_06086_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14087_ (.A1(_04645_),
    .A2(_06086_),
    .A3(_05992_),
    .ZN(_06087_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14088_ (.A1(_05440_),
    .A2(_05980_),
    .A3(_05994_),
    .ZN(_06088_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _14089_ (.A1(_06087_),
    .A2(_06088_),
    .Z(_06089_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14090_ (.A1(_06002_),
    .A2(_06021_),
    .ZN(_06090_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _14091_ (.A1(_06004_),
    .A2(_06020_),
    .B(_06090_),
    .ZN(_06091_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14092_ (.A1(_04561_),
    .A2(_06086_),
    .ZN(_06092_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14093_ (.I(_06005_),
    .Z(_06093_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14094_ (.A1(_05446_),
    .A2(_06093_),
    .A3(_06010_),
    .ZN(_06094_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _14095_ (.A1(_06007_),
    .A2(_06009_),
    .B(_06094_),
    .ZN(_06095_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14096_ (.I(_06005_),
    .Z(_06096_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14097_ (.A1(_04416_),
    .A2(_06096_),
    .ZN(_06097_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _14098_ (.A1(_06095_),
    .A2(_06097_),
    .ZN(_06098_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14099_ (.A1(_06092_),
    .A2(_06098_),
    .Z(_06099_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _14100_ (.A1(_06091_),
    .A2(_06099_),
    .ZN(_06100_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14101_ (.A1(_06089_),
    .A2(_06100_),
    .Z(_06101_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14102_ (.A1(_06024_),
    .A2(_06055_),
    .ZN(_06102_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _14103_ (.A1(_06022_),
    .A2(_06056_),
    .B(_06102_),
    .ZN(_06103_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _14104_ (.A1(_06026_),
    .A2(_06041_),
    .Z(_06104_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _14105_ (.A1(_06042_),
    .A2(_06054_),
    .B(_06104_),
    .ZN(_06105_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14106_ (.A1(_06030_),
    .A2(_06035_),
    .ZN(_06106_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _14107_ (.A1(_06036_),
    .A2(_06040_),
    .B(_06106_),
    .ZN(_06107_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _14108_ (.A1(_06031_),
    .A2(_06032_),
    .Z(_06108_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _14109_ (.A1(_06033_),
    .A2(_06034_),
    .B(_06108_),
    .ZN(_06109_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14110_ (.A1(_03397_),
    .A2(_04402_),
    .A3(_05106_),
    .ZN(_06110_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14111_ (.A1(_03413_),
    .A2(_04488_),
    .A3(net58),
    .ZN(_06111_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _14112_ (.A1(_06110_),
    .A2(_06111_),
    .ZN(_06112_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14113_ (.A1(_04711_),
    .A2(_04817_),
    .ZN(_06113_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _14114_ (.A1(_06112_),
    .A2(_06113_),
    .ZN(_06114_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _14115_ (.A1(_06109_),
    .A2(_06114_),
    .ZN(_06115_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14116_ (.A1(_04740_),
    .A2(_04781_),
    .ZN(_06116_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14117_ (.A1(_04803_),
    .A2(_04861_),
    .ZN(_06117_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _14118_ (.A1(_06116_),
    .A2(_06117_),
    .ZN(_06118_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _14119_ (.A1(_04801_),
    .A2(_04927_),
    .ZN(_06119_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14120_ (.A1(_06118_),
    .A2(_06119_),
    .Z(_06120_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14121_ (.A1(_06115_),
    .A2(_06120_),
    .Z(_06121_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14122_ (.A1(_06107_),
    .A2(_06121_),
    .Z(_06122_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _14123_ (.A1(_06049_),
    .A2(_06050_),
    .Z(_06123_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _14124_ (.A1(_06049_),
    .A2(_06050_),
    .Z(_06124_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _14125_ (.A1(_06123_),
    .A2(_06051_),
    .B(_06124_),
    .ZN(_06125_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _14126_ (.A1(_06038_),
    .A2(_06039_),
    .Z(_06126_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _14127_ (.A1(_06038_),
    .A2(_06039_),
    .Z(_06127_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _14128_ (.A1(_06037_),
    .A2(_06126_),
    .B(_06127_),
    .ZN(_06128_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14129_ (.A1(_04376_),
    .A2(_05077_),
    .ZN(_06129_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14130_ (.A1(_04371_),
    .A2(_05185_),
    .ZN(_06130_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14131_ (.A1(_04367_),
    .A2(_05347_),
    .ZN(_06131_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _14132_ (.A1(_06129_),
    .A2(_06130_),
    .A3(_06131_),
    .ZN(_06132_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14133_ (.A1(_06128_),
    .A2(_06132_),
    .Z(_06133_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14134_ (.A1(_06125_),
    .A2(_06133_),
    .Z(_06134_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _14135_ (.A1(_06122_),
    .A2(_06134_),
    .ZN(_06135_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _14136_ (.A1(_06105_),
    .A2(_06135_),
    .ZN(_06136_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14137_ (.A1(_06014_),
    .A2(_06018_),
    .ZN(_06137_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14138_ (.A1(_06011_),
    .A2(_06019_),
    .ZN(_06138_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14139_ (.A1(_06137_),
    .A2(_06138_),
    .ZN(_06139_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _14140_ (.I(_06052_),
    .ZN(_06140_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14141_ (.A1(_06045_),
    .A2(_06053_),
    .ZN(_06141_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _14142_ (.A1(_06048_),
    .A2(_06140_),
    .B(_06141_),
    .ZN(_06142_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14143_ (.A1(_04529_),
    .A2(_06008_),
    .ZN(_06143_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14144_ (.A1(_04742_),
    .A2(_05690_),
    .ZN(_06144_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14145_ (.A1(\filters.band[26] ),
    .A2(_04186_),
    .ZN(_06145_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14146_ (.A1(_06144_),
    .A2(_06145_),
    .Z(_06146_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _14147_ (.A1(_06143_),
    .A2(_06146_),
    .ZN(_06147_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _14148_ (.A1(_06015_),
    .A2(_06016_),
    .Z(_06148_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _14149_ (.A1(_06015_),
    .A2(_06016_),
    .Z(_06149_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _14150_ (.A1(_06148_),
    .A2(_06017_),
    .B(_06149_),
    .ZN(_06150_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14151_ (.A1(_05069_),
    .A2(_05350_),
    .ZN(_06151_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14152_ (.A1(_04258_),
    .A2(_05504_),
    .ZN(_06152_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14153_ (.A1(_06151_),
    .A2(_06152_),
    .Z(_06153_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14154_ (.A1(_04230_),
    .A2(_05588_),
    .ZN(_06154_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _14155_ (.A1(_06153_),
    .A2(_06154_),
    .ZN(_06155_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14156_ (.A1(_06150_),
    .A2(_06155_),
    .Z(_06156_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _14157_ (.A1(_06147_),
    .A2(_06156_),
    .ZN(_06157_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14158_ (.A1(_06142_),
    .A2(_06157_),
    .Z(_06158_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _14159_ (.A1(_06139_),
    .A2(_06158_),
    .ZN(_06159_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14160_ (.A1(_06136_),
    .A2(_06159_),
    .Z(_06160_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14161_ (.A1(_06103_),
    .A2(_06160_),
    .Z(_06161_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _14162_ (.A1(_06101_),
    .A2(_06161_),
    .ZN(_06162_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _14163_ (.A1(_06085_),
    .A2(_06162_),
    .Z(_06163_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _14164_ (.A1(_06082_),
    .A2(_06163_),
    .ZN(_06164_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14165_ (.A1(_05979_),
    .A2(_06058_),
    .ZN(_06165_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14166_ (.A1(_05979_),
    .A2(_06058_),
    .ZN(_06166_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _14167_ (.A1(_05977_),
    .A2(_06165_),
    .B(_06166_),
    .ZN(_06167_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _14168_ (.A1(_06164_),
    .A2(_06167_),
    .Z(_06168_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14169_ (.A1(_05967_),
    .A2(_06062_),
    .ZN(_06169_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _14170_ (.I(_06169_),
    .ZN(_06170_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14171_ (.A1(_06059_),
    .A2(_06061_),
    .ZN(_06171_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14172_ (.A1(_06059_),
    .A2(_06061_),
    .ZN(_06172_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _14173_ (.A1(_06063_),
    .A2(_06171_),
    .B(_06172_),
    .ZN(_06173_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _14174_ (.I(_06173_),
    .ZN(_06174_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _14175_ (.A1(_05877_),
    .A2(_06170_),
    .B(_06174_),
    .ZN(_06175_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14176_ (.A1(_06168_),
    .A2(_06175_),
    .Z(_06176_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _14177_ (.I(_06066_),
    .Z(_06177_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14178_ (.A1(_03329_),
    .A2(_05853_),
    .ZN(_06178_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _14179_ (.A1(_03330_),
    .A2(_06177_),
    .B(_06178_),
    .ZN(_06179_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14180_ (.A1(_06176_),
    .A2(_06179_),
    .Z(_06180_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _14181_ (.I(_06070_),
    .ZN(_06181_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _14182_ (.A1(_05972_),
    .A2(_06070_),
    .A3(_06071_),
    .ZN(_06182_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _14183_ (.A1(_06074_),
    .A2(_06181_),
    .B1(_06182_),
    .B2(_05869_),
    .C(_06071_),
    .ZN(_06183_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _14184_ (.A1(_06180_),
    .A2(_06183_),
    .ZN(_06184_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14185_ (.A1(_05975_),
    .A2(_06184_),
    .ZN(_06185_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _14186_ (.I(_01821_),
    .Z(_06186_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _14187_ (.I(_06186_),
    .Z(_06187_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _14188_ (.A1(_03330_),
    .A2(_06080_),
    .B(_06185_),
    .C(_06187_),
    .ZN(_00532_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _14189_ (.A1(_06091_),
    .A2(_06099_),
    .Z(_06188_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _14190_ (.A1(_06089_),
    .A2(_06100_),
    .B(_06188_),
    .ZN(_06189_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14191_ (.A1(_06103_),
    .A2(_06160_),
    .ZN(_06190_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14192_ (.A1(_06101_),
    .A2(_06161_),
    .ZN(_06191_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14193_ (.A1(_06190_),
    .A2(_06191_),
    .ZN(_06192_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _14194_ (.A1(_06105_),
    .A2(_06135_),
    .Z(_06193_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _14195_ (.A1(_06136_),
    .A2(_06159_),
    .B(_06193_),
    .ZN(_06194_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14196_ (.A1(_06107_),
    .A2(_06121_),
    .ZN(_06195_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14197_ (.A1(_06122_),
    .A2(_06134_),
    .ZN(_06196_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _14198_ (.A1(_06195_),
    .A2(_06196_),
    .ZN(_06197_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _14199_ (.I(_06114_),
    .ZN(_06198_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14200_ (.A1(_06109_),
    .A2(_06198_),
    .ZN(_06199_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14201_ (.A1(_06115_),
    .A2(_06120_),
    .ZN(_06200_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14202_ (.A1(_06199_),
    .A2(_06200_),
    .ZN(_06201_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14203_ (.A1(_06110_),
    .A2(_06111_),
    .ZN(_06202_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14204_ (.A1(_06112_),
    .A2(_06113_),
    .ZN(_06203_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _14205_ (.A1(_06202_),
    .A2(_06203_),
    .ZN(_06204_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14206_ (.A1(_04750_),
    .A2(_05625_),
    .ZN(_06205_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14207_ (.A1(_04737_),
    .A2(_05731_),
    .ZN(_06206_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _14208_ (.A1(_06205_),
    .A2(_06206_),
    .ZN(_06207_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14209_ (.A1(_05183_),
    .A2(_04819_),
    .ZN(_06208_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _14210_ (.A1(_06207_),
    .A2(_06208_),
    .ZN(_06209_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _14211_ (.A1(_06204_),
    .A2(_06209_),
    .ZN(_06210_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _14212_ (.A1(_05465_),
    .A2(_05049_),
    .ZN(_06211_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14213_ (.A1(_05930_),
    .A2(_05075_),
    .ZN(_06212_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _14214_ (.A1(_04896_),
    .A2(_05181_),
    .ZN(_06213_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _14215_ (.A1(_06211_),
    .A2(_06212_),
    .A3(_06213_),
    .ZN(_06214_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14216_ (.A1(_06210_),
    .A2(_06214_),
    .Z(_06215_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14217_ (.A1(_06201_),
    .A2(_06215_),
    .Z(_06216_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _14218_ (.A1(_06129_),
    .A2(_06130_),
    .Z(_06217_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _14219_ (.A1(_06129_),
    .A2(_06130_),
    .Z(_06218_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _14220_ (.A1(_06217_),
    .A2(_06131_),
    .B(_06218_),
    .ZN(_06219_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _14221_ (.A1(_06116_),
    .A2(_06117_),
    .Z(_06220_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _14222_ (.A1(_06118_),
    .A2(_06119_),
    .B(_06220_),
    .ZN(_06221_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14223_ (.A1(_04326_),
    .A2(_05501_),
    .ZN(_06222_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14224_ (.A1(_04452_),
    .A2(_05947_),
    .ZN(_06223_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14225_ (.A1(_04893_),
    .A2(_05447_),
    .ZN(_06224_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14226_ (.A1(_06223_),
    .A2(_06224_),
    .Z(_06225_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _14227_ (.A1(_06222_),
    .A2(_06225_),
    .ZN(_06226_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14228_ (.A1(_06221_),
    .A2(_06226_),
    .Z(_06227_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14229_ (.A1(_06219_),
    .A2(_06227_),
    .Z(_06228_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14230_ (.A1(_06216_),
    .A2(_06228_),
    .Z(_06229_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14231_ (.A1(_06197_),
    .A2(_06229_),
    .Z(_06230_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14232_ (.A1(_06150_),
    .A2(_06155_),
    .ZN(_06231_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14233_ (.A1(_06147_),
    .A2(_06156_),
    .ZN(_06232_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14234_ (.A1(_06231_),
    .A2(_06232_),
    .ZN(_06233_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14235_ (.A1(_06128_),
    .A2(_06132_),
    .ZN(_06234_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14236_ (.A1(_06125_),
    .A2(_06133_),
    .ZN(_06235_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14237_ (.A1(_06234_),
    .A2(_06235_),
    .ZN(_06236_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14238_ (.A1(\filters.band[26] ),
    .A2(_04596_),
    .ZN(_06237_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14239_ (.A1(_04504_),
    .A2(_05989_),
    .ZN(_06238_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14240_ (.A1(\filters.band[27] ),
    .A2(_04599_),
    .ZN(_06239_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _14241_ (.A1(_06237_),
    .A2(_06238_),
    .A3(_06239_),
    .ZN(_06240_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14242_ (.A1(_04575_),
    .A2(_05774_),
    .A3(_06153_),
    .ZN(_06241_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _14243_ (.A1(_06151_),
    .A2(_06152_),
    .B(_06241_),
    .ZN(_06242_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14244_ (.A1(_04699_),
    .A2(_05505_),
    .ZN(_06243_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14245_ (.A1(_04697_),
    .A2(_05687_),
    .ZN(_06244_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14246_ (.A1(_06243_),
    .A2(_06244_),
    .Z(_06245_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14247_ (.A1(_04231_),
    .A2(_05891_),
    .ZN(_06246_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _14248_ (.A1(_06245_),
    .A2(_06246_),
    .ZN(_06247_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14249_ (.A1(_06242_),
    .A2(_06247_),
    .Z(_06248_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14250_ (.A1(_06240_),
    .A2(_06248_),
    .Z(_06249_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14251_ (.A1(_06236_),
    .A2(_06249_),
    .Z(_06250_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14252_ (.A1(_06233_),
    .A2(_06250_),
    .Z(_06251_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14253_ (.A1(_06230_),
    .A2(_06251_),
    .Z(_06252_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14254_ (.A1(_06194_),
    .A2(_06252_),
    .Z(_06253_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14255_ (.I(_05560_),
    .Z(_06254_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14256_ (.A1(_06254_),
    .A2(_06096_),
    .A3(_06095_),
    .ZN(_06255_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14257_ (.A1(_05982_),
    .A2(_06086_),
    .A3(_06098_),
    .ZN(_06256_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _14258_ (.A1(_06255_),
    .A2(_06256_),
    .Z(_06257_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14259_ (.A1(_06142_),
    .A2(_06157_),
    .ZN(_06258_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _14260_ (.A1(_06139_),
    .A2(_06158_),
    .B(_06258_),
    .ZN(_06259_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _14261_ (.A1(_06144_),
    .A2(_06145_),
    .Z(_06260_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14262_ (.I(_06008_),
    .Z(_06261_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14263_ (.A1(_04616_),
    .A2(_06261_),
    .A3(_06146_),
    .ZN(_06262_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _14264_ (.A1(_06260_),
    .A2(_06262_),
    .Z(_06263_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14265_ (.A1(_04644_),
    .A2(_06261_),
    .ZN(_06264_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _14266_ (.A1(_06263_),
    .A2(_06264_),
    .ZN(_06265_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14267_ (.A1(_05440_),
    .A2(_06096_),
    .ZN(_06266_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _14268_ (.A1(_06265_),
    .A2(_06266_),
    .Z(_06267_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14269_ (.A1(_06265_),
    .A2(_06266_),
    .ZN(_06268_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14270_ (.A1(_06267_),
    .A2(_06268_),
    .ZN(_06269_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _14271_ (.A1(_06259_),
    .A2(_06269_),
    .Z(_06270_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14272_ (.A1(_06259_),
    .A2(_06269_),
    .ZN(_06271_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14273_ (.A1(_06270_),
    .A2(_06271_),
    .ZN(_06272_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14274_ (.A1(_06257_),
    .A2(_06272_),
    .Z(_06273_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14275_ (.A1(_06253_),
    .A2(_06273_),
    .Z(_06274_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _14276_ (.A1(_06189_),
    .A2(_06192_),
    .A3(_06274_),
    .ZN(_06275_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14277_ (.A1(_06085_),
    .A2(_06162_),
    .ZN(_06276_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _14278_ (.A1(_06082_),
    .A2(_06163_),
    .B(_06276_),
    .ZN(_06277_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14279_ (.A1(_06275_),
    .A2(_06277_),
    .Z(_06278_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _14280_ (.I(_06168_),
    .ZN(_06279_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14281_ (.A1(_06164_),
    .A2(_06167_),
    .ZN(_06280_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _14282_ (.I(_06280_),
    .ZN(_06281_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _14283_ (.A1(_06279_),
    .A2(_06175_),
    .B(_06281_),
    .ZN(_06282_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _14284_ (.A1(_06278_),
    .A2(_06282_),
    .ZN(_06283_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14285_ (.A1(_03345_),
    .A2(_05853_),
    .ZN(_06284_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _14286_ (.A1(_03347_),
    .A2(_06177_),
    .B(_06284_),
    .ZN(_06285_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14287_ (.A1(_06283_),
    .A2(_06285_),
    .Z(_06286_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14288_ (.I(_06176_),
    .Z(_06287_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14289_ (.A1(_06287_),
    .A2(_06179_),
    .ZN(_06288_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14290_ (.A1(_06287_),
    .A2(_06179_),
    .ZN(_06289_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _14291_ (.A1(_06288_),
    .A2(_06183_),
    .B(_06289_),
    .ZN(_06290_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14292_ (.A1(_06286_),
    .A2(_06290_),
    .Z(_06291_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14293_ (.A1(_05975_),
    .A2(_06291_),
    .ZN(_06292_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _14294_ (.A1(_03347_),
    .A2(_06080_),
    .B(_06292_),
    .C(_06187_),
    .ZN(_00533_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _14295_ (.I(_06283_),
    .Z(_06293_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _14296_ (.I(_06293_),
    .Z(_06294_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14297_ (.A1(_06294_),
    .A2(_06285_),
    .ZN(_06295_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _14298_ (.A1(_06287_),
    .A2(_06179_),
    .B1(_06293_),
    .B2(_06285_),
    .ZN(_06296_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14299_ (.A1(_06180_),
    .A2(_06286_),
    .ZN(_06297_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_4 _14300_ (.A1(_06295_),
    .A2(_06296_),
    .B1(_06297_),
    .B2(_06183_),
    .ZN(_06298_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14301_ (.A1(_06168_),
    .A2(_06278_),
    .ZN(_06299_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _14302_ (.A1(_06169_),
    .A2(_06299_),
    .ZN(_06300_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _14303_ (.A1(_06275_),
    .A2(_06277_),
    .Z(_06301_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _14304_ (.A1(_06281_),
    .A2(_06301_),
    .B1(_06299_),
    .B2(_06173_),
    .ZN(_06302_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14305_ (.A1(_06275_),
    .A2(_06277_),
    .ZN(_06303_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _14306_ (.A1(_05877_),
    .A2(_06300_),
    .B(_06302_),
    .C(_06303_),
    .ZN(_06304_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _14307_ (.A1(_06257_),
    .A2(_06272_),
    .B(_06270_),
    .ZN(_06305_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14308_ (.A1(_06194_),
    .A2(_06252_),
    .ZN(_06306_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14309_ (.A1(_06253_),
    .A2(_06273_),
    .ZN(_06307_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14310_ (.A1(_06306_),
    .A2(_06307_),
    .ZN(_06308_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14311_ (.A1(_06197_),
    .A2(_06229_),
    .ZN(_06309_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14312_ (.A1(_06230_),
    .A2(_06251_),
    .ZN(_06310_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14313_ (.A1(_06309_),
    .A2(_06310_),
    .ZN(_06311_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14314_ (.A1(_06201_),
    .A2(_06215_),
    .ZN(_06312_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14315_ (.A1(_06216_),
    .A2(_06228_),
    .ZN(_06313_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14316_ (.A1(_06312_),
    .A2(_06313_),
    .ZN(_06314_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _14317_ (.A1(_06210_),
    .A2(_06214_),
    .Z(_06315_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _14318_ (.A1(_06204_),
    .A2(_06209_),
    .B(_06315_),
    .ZN(_06316_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14319_ (.A1(_06205_),
    .A2(_06206_),
    .ZN(_06317_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14320_ (.A1(_06207_),
    .A2(_06208_),
    .ZN(_06318_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14321_ (.A1(_06317_),
    .A2(_06318_),
    .ZN(_06319_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14322_ (.A1(_05469_),
    .A2(_06027_),
    .ZN(_06320_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14323_ (.A1(_04858_),
    .A2(_05487_),
    .ZN(_06321_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _14324_ (.A1(_06320_),
    .A2(_06321_),
    .ZN(_06322_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14325_ (.A1(_04820_),
    .A2(_04924_),
    .ZN(_06323_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _14326_ (.A1(_06322_),
    .A2(_06323_),
    .ZN(_06324_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _14327_ (.A1(_06319_),
    .A2(_06324_),
    .ZN(_06325_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14328_ (.A1(_05909_),
    .A2(_05092_),
    .ZN(_06326_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14329_ (.A1(_04806_),
    .A2(_05280_),
    .ZN(_06327_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14330_ (.A1(_04446_),
    .A2(_05367_),
    .ZN(_06328_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _14331_ (.A1(_06326_),
    .A2(_06327_),
    .A3(_06328_),
    .Z(_06329_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14332_ (.A1(_06325_),
    .A2(_06329_),
    .Z(_06330_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14333_ (.A1(_06316_),
    .A2(_06330_),
    .Z(_06331_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14334_ (.I(_04355_),
    .Z(_06332_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14335_ (.A1(_06332_),
    .A2(_05570_),
    .A3(_06225_),
    .ZN(_06333_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _14336_ (.A1(_06223_),
    .A2(_06224_),
    .B(_06333_),
    .ZN(_06334_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14337_ (.A1(_06211_),
    .A2(_06212_),
    .ZN(_06335_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14338_ (.A1(_06211_),
    .A2(_06212_),
    .ZN(_06336_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _14339_ (.A1(_06335_),
    .A2(_06213_),
    .B(_06336_),
    .ZN(_06337_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14340_ (.A1(_04326_),
    .A2(_05585_),
    .ZN(_06338_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14341_ (.A1(_04378_),
    .A2(_05447_),
    .ZN(_06339_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14342_ (.A1(_04318_),
    .A2(_05500_),
    .ZN(_06340_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14343_ (.A1(_06339_),
    .A2(_06340_),
    .Z(_06341_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _14344_ (.A1(_06338_),
    .A2(_06341_),
    .ZN(_06342_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14345_ (.A1(_06337_),
    .A2(_06342_),
    .Z(_06343_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _14346_ (.I(_06343_),
    .ZN(_06344_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14347_ (.A1(_06334_),
    .A2(_06344_),
    .Z(_06345_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14348_ (.A1(_06331_),
    .A2(_06345_),
    .Z(_06346_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14349_ (.A1(_06314_),
    .A2(_06346_),
    .Z(_06347_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14350_ (.A1(_06242_),
    .A2(_06247_),
    .ZN(_06348_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14351_ (.A1(_06240_),
    .A2(_06248_),
    .ZN(_06349_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14352_ (.A1(_06348_),
    .A2(_06349_),
    .ZN(_06350_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14353_ (.A1(_06221_),
    .A2(_06226_),
    .ZN(_06351_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14354_ (.A1(_06219_),
    .A2(_06227_),
    .ZN(_06352_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14355_ (.A1(_06351_),
    .A2(_06352_),
    .ZN(_06353_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14356_ (.A1(\filters.band[27] ),
    .A2(_04578_),
    .ZN(_06354_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14357_ (.A1(_04600_),
    .A2(_06093_),
    .ZN(_06355_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14358_ (.I(\filters.band[28] ),
    .Z(_06356_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14359_ (.A1(_06356_),
    .A2(_04617_),
    .ZN(_06357_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _14360_ (.A1(_06354_),
    .A2(_06355_),
    .A3(_06357_),
    .ZN(_06358_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14361_ (.I(_04575_),
    .Z(_06359_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14362_ (.A1(_06359_),
    .A2(_05891_),
    .A3(_06245_),
    .ZN(_06360_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _14363_ (.A1(_06243_),
    .A2(_06244_),
    .B(_06360_),
    .ZN(_06361_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14364_ (.A1(_06359_),
    .A2(_05989_),
    .ZN(_06362_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14365_ (.A1(_05509_),
    .A2(_05774_),
    .ZN(_06363_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14366_ (.A1(_04222_),
    .A2(_05793_),
    .ZN(_06364_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14367_ (.A1(_06363_),
    .A2(_06364_),
    .Z(_06365_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _14368_ (.A1(_06362_),
    .A2(_06365_),
    .ZN(_06366_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14369_ (.A1(_06361_),
    .A2(_06366_),
    .Z(_06367_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14370_ (.A1(_06358_),
    .A2(_06367_),
    .Z(_06368_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14371_ (.A1(_06353_),
    .A2(_06368_),
    .Z(_06369_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14372_ (.A1(_06350_),
    .A2(_06369_),
    .Z(_06370_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14373_ (.A1(_06347_),
    .A2(_06370_),
    .Z(_06371_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14374_ (.A1(_06311_),
    .A2(_06371_),
    .Z(_06372_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _14375_ (.A1(_06263_),
    .A2(_06264_),
    .B(_06267_),
    .ZN(_06373_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14376_ (.A1(_06236_),
    .A2(_06249_),
    .ZN(_06374_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14377_ (.A1(_06233_),
    .A2(_06250_),
    .ZN(_06375_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14378_ (.A1(_06374_),
    .A2(_06375_),
    .ZN(_06376_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _14379_ (.A1(_06238_),
    .A2(_06239_),
    .Z(_06377_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _14380_ (.A1(_06238_),
    .A2(_06239_),
    .Z(_06378_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _14381_ (.A1(_06237_),
    .A2(_06377_),
    .B(_06378_),
    .ZN(_06379_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _14382_ (.I(\filters.band[26] ),
    .Z(_06380_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14383_ (.A1(_06380_),
    .A2(_04632_),
    .ZN(_06381_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _14384_ (.A1(_06379_),
    .A2(_06381_),
    .ZN(_06382_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14385_ (.I(_06261_),
    .Z(_06383_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14386_ (.A1(_05563_),
    .A2(_06383_),
    .ZN(_06384_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _14387_ (.A1(_06382_),
    .A2(_06384_),
    .ZN(_06385_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14388_ (.A1(_06376_),
    .A2(_06385_),
    .Z(_06386_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14389_ (.A1(_06373_),
    .A2(_06386_),
    .Z(_06387_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14390_ (.A1(_06372_),
    .A2(_06387_),
    .Z(_06388_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14391_ (.A1(_06308_),
    .A2(_06388_),
    .Z(_06389_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14392_ (.A1(_06305_),
    .A2(_06389_),
    .Z(_06390_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14393_ (.A1(_06192_),
    .A2(_06274_),
    .ZN(_06391_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _14394_ (.A1(_06192_),
    .A2(_06274_),
    .Z(_06392_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14395_ (.A1(_06189_),
    .A2(_06391_),
    .A3(_06392_),
    .ZN(_06393_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14396_ (.A1(_06391_),
    .A2(_06393_),
    .ZN(_06394_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _14397_ (.A1(_06390_),
    .A2(_06394_),
    .ZN(_06395_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _14398_ (.A1(net51),
    .A2(_06395_),
    .ZN(_06396_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _14399_ (.I(_05853_),
    .Z(_06397_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14400_ (.A1(_03360_),
    .A2(_03221_),
    .ZN(_06398_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _14401_ (.A1(_03361_),
    .A2(_06397_),
    .B(_06398_),
    .ZN(_06399_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14402_ (.A1(_06396_),
    .A2(_06399_),
    .Z(_06400_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14403_ (.A1(_06298_),
    .A2(_06400_),
    .Z(_06401_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14404_ (.A1(_05975_),
    .A2(_06401_),
    .ZN(_06402_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _14405_ (.A1(_03361_),
    .A2(_06080_),
    .B(_06402_),
    .C(_06187_),
    .ZN(_00534_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14406_ (.I(_05543_),
    .Z(_06403_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14407_ (.A1(_06376_),
    .A2(_06385_),
    .ZN(_06404_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14408_ (.A1(_06373_),
    .A2(_06386_),
    .ZN(_06405_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14409_ (.A1(_06404_),
    .A2(_06405_),
    .ZN(_06406_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14410_ (.A1(_06311_),
    .A2(_06371_),
    .ZN(_06407_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14411_ (.A1(_06372_),
    .A2(_06387_),
    .ZN(_06408_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14412_ (.A1(_06407_),
    .A2(_06408_),
    .ZN(_06409_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14413_ (.A1(_06314_),
    .A2(_06346_),
    .ZN(_06410_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14414_ (.A1(_06347_),
    .A2(_06370_),
    .ZN(_06411_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14415_ (.A1(_06410_),
    .A2(_06411_),
    .ZN(_06412_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14416_ (.A1(_06316_),
    .A2(_06330_),
    .ZN(_06413_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14417_ (.A1(_06331_),
    .A2(_06345_),
    .ZN(_06414_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14418_ (.A1(_06413_),
    .A2(_06414_),
    .ZN(_06415_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _14419_ (.A1(_06319_),
    .A2(_06324_),
    .Z(_06416_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _14420_ (.A1(_06325_),
    .A2(_06329_),
    .B(_06416_),
    .ZN(_06417_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14421_ (.A1(_06320_),
    .A2(_06321_),
    .ZN(_06418_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14422_ (.A1(_06322_),
    .A2(_06323_),
    .ZN(_06419_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _14423_ (.A1(_06418_),
    .A2(_06419_),
    .ZN(_06420_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14424_ (.A1(_05183_),
    .A2(_06027_),
    .ZN(_06421_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14425_ (.A1(_04923_),
    .A2(_05732_),
    .ZN(_06422_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14426_ (.A1(_04819_),
    .A2(_05075_),
    .ZN(_06423_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _14427_ (.A1(_06421_),
    .A2(_06422_),
    .A3(_06423_),
    .Z(_06424_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14428_ (.A1(_06420_),
    .A2(_06424_),
    .Z(_06425_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14429_ (.A1(_05721_),
    .A2(_05079_),
    .ZN(_06426_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14430_ (.A1(_04805_),
    .A2(_05187_),
    .ZN(_06427_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14431_ (.A1(_06426_),
    .A2(_06427_),
    .Z(_06428_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14432_ (.A1(_04802_),
    .A2(_05448_),
    .ZN(_06429_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _14433_ (.A1(_06428_),
    .A2(_06429_),
    .ZN(_06430_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14434_ (.A1(_06425_),
    .A2(_06430_),
    .Z(_06431_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14435_ (.A1(_06417_),
    .A2(_06431_),
    .Z(_06432_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _14436_ (.A1(_06339_),
    .A2(_06340_),
    .Z(_06433_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14437_ (.A1(_06332_),
    .A2(_05671_),
    .A3(_06341_),
    .ZN(_06434_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _14438_ (.A1(_06433_),
    .A2(_06434_),
    .Z(_06435_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _14439_ (.A1(_06326_),
    .A2(_06327_),
    .Z(_06436_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _14440_ (.A1(_06326_),
    .A2(_06327_),
    .Z(_06437_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _14441_ (.A1(_06436_),
    .A2(_06328_),
    .B(_06437_),
    .ZN(_06438_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14442_ (.A1(_04355_),
    .A2(_05774_),
    .ZN(_06439_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14443_ (.A1(_04453_),
    .A2(_05500_),
    .ZN(_06440_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14444_ (.A1(_04318_),
    .A2(_05585_),
    .ZN(_06441_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14445_ (.A1(_06440_),
    .A2(_06441_),
    .Z(_06442_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _14446_ (.A1(_06439_),
    .A2(_06442_),
    .ZN(_06443_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _14447_ (.A1(_06438_),
    .A2(_06443_),
    .ZN(_06444_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14448_ (.A1(_06435_),
    .A2(_06444_),
    .Z(_06445_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14449_ (.A1(_06432_),
    .A2(_06445_),
    .Z(_06446_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14450_ (.A1(_06415_),
    .A2(_06446_),
    .Z(_06447_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14451_ (.A1(_06361_),
    .A2(_06366_),
    .ZN(_06448_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14452_ (.A1(_06358_),
    .A2(_06367_),
    .ZN(_06449_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14453_ (.A1(_06448_),
    .A2(_06449_),
    .ZN(_06450_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _14454_ (.I(_06342_),
    .ZN(_06451_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14455_ (.A1(_06334_),
    .A2(_06344_),
    .ZN(_06452_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _14456_ (.A1(_06337_),
    .A2(_06451_),
    .B(_06452_),
    .ZN(_06453_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14457_ (.A1(\filters.band[28] ),
    .A2(_05446_),
    .ZN(_06454_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14458_ (.A1(_04600_),
    .A2(_06261_),
    .ZN(_06455_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _14459_ (.I(\filters.band[29] ),
    .Z(_06456_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14460_ (.A1(_06456_),
    .A2(_04617_),
    .ZN(_06457_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _14461_ (.A1(_06454_),
    .A2(_06455_),
    .A3(_06457_),
    .ZN(_06458_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14462_ (.A1(_04576_),
    .A2(_05990_),
    .A3(_06365_),
    .ZN(_06459_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _14463_ (.A1(_06363_),
    .A2(_06364_),
    .B(_06459_),
    .ZN(_06460_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14464_ (.A1(_06359_),
    .A2(_06093_),
    .ZN(_06461_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14465_ (.A1(_05509_),
    .A2(_05793_),
    .ZN(_06462_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14466_ (.A1(_05510_),
    .A2(_05989_),
    .ZN(_06463_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14467_ (.A1(_06462_),
    .A2(_06463_),
    .Z(_06464_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _14468_ (.A1(_06461_),
    .A2(_06464_),
    .ZN(_06465_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14469_ (.A1(_06460_),
    .A2(_06465_),
    .Z(_06466_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14470_ (.A1(_06458_),
    .A2(_06466_),
    .Z(_06467_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14471_ (.A1(_06453_),
    .A2(_06467_),
    .Z(_06468_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14472_ (.A1(_06450_),
    .A2(_06468_),
    .Z(_06469_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14473_ (.A1(_06447_),
    .A2(_06469_),
    .Z(_06470_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14474_ (.A1(_06412_),
    .A2(_06470_),
    .Z(_06471_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _14475_ (.I(_06380_),
    .Z(_06472_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14476_ (.I(_06254_),
    .Z(_06473_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14477_ (.A1(_06472_),
    .A2(_06473_),
    .A3(_06379_),
    .ZN(_06474_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14478_ (.A1(_05982_),
    .A2(_06383_),
    .A3(_06382_),
    .ZN(_06475_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _14479_ (.A1(_06474_),
    .A2(_06475_),
    .Z(_06476_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14480_ (.A1(_06353_),
    .A2(_06368_),
    .ZN(_06477_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14481_ (.A1(_06350_),
    .A2(_06369_),
    .ZN(_06478_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14482_ (.A1(_06477_),
    .A2(_06478_),
    .ZN(_06479_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14483_ (.A1(_06380_),
    .A2(_05563_),
    .ZN(_06480_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _14484_ (.A1(_06355_),
    .A2(_06357_),
    .Z(_06481_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _14485_ (.A1(_06355_),
    .A2(_06357_),
    .Z(_06482_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _14486_ (.A1(_06354_),
    .A2(_06481_),
    .B(_06482_),
    .ZN(_06483_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _14487_ (.I(\filters.band[27] ),
    .Z(_06484_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14488_ (.A1(_06484_),
    .A2(_05560_),
    .ZN(_06485_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _14489_ (.A1(_06480_),
    .A2(_06483_),
    .A3(_06485_),
    .Z(_06486_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _14490_ (.A1(_06479_),
    .A2(_06486_),
    .ZN(_06487_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14491_ (.A1(_06476_),
    .A2(_06487_),
    .Z(_06488_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14492_ (.A1(_06471_),
    .A2(_06488_),
    .Z(_06489_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _14493_ (.A1(_06406_),
    .A2(_06409_),
    .A3(_06489_),
    .ZN(_06490_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14494_ (.A1(_06308_),
    .A2(_06388_),
    .ZN(_06491_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14495_ (.A1(_06305_),
    .A2(_06389_),
    .ZN(_06492_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14496_ (.A1(_06491_),
    .A2(_06492_),
    .ZN(_06493_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14497_ (.A1(_06490_),
    .A2(_06493_),
    .Z(_06494_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _14498_ (.A1(_06390_),
    .A2(_06394_),
    .Z(_06495_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _14499_ (.I(_06495_),
    .ZN(_06496_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _14500_ (.A1(_06304_),
    .A2(_06395_),
    .B(_06496_),
    .ZN(_06497_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14501_ (.A1(_06494_),
    .A2(_06497_),
    .Z(_06498_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _14502_ (.I(_06498_),
    .Z(_06499_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14503_ (.A1(_03374_),
    .A2(_06177_),
    .ZN(_06500_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _14504_ (.A1(_03380_),
    .A2(_03378_),
    .B(_06500_),
    .ZN(_06501_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14505_ (.A1(_06499_),
    .A2(_06501_),
    .Z(_06502_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14506_ (.A1(_06396_),
    .A2(_06399_),
    .ZN(_06503_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14507_ (.A1(_06298_),
    .A2(_06400_),
    .ZN(_06504_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14508_ (.A1(_06503_),
    .A2(_06504_),
    .ZN(_06505_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14509_ (.A1(_06502_),
    .A2(_06505_),
    .Z(_06506_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14510_ (.A1(_06403_),
    .A2(_06506_),
    .ZN(_06507_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _14511_ (.A1(_03380_),
    .A2(_06080_),
    .B(_06507_),
    .C(_06187_),
    .ZN(_00535_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _14512_ (.I(_05544_),
    .Z(_06508_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _14513_ (.A1(_06491_),
    .A2(_06492_),
    .B(_06490_),
    .ZN(_06509_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14514_ (.A1(_06491_),
    .A2(_06492_),
    .A3(_06490_),
    .ZN(_06510_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _14515_ (.A1(_06495_),
    .A2(_06509_),
    .B(_06510_),
    .ZN(_06511_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _14516_ (.A1(_06304_),
    .A2(_06395_),
    .A3(_06494_),
    .B(_06511_),
    .ZN(_06512_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _14517_ (.A1(_06409_),
    .A2(_06489_),
    .Z(_06513_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _14518_ (.A1(_06409_),
    .A2(_06489_),
    .Z(_06514_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _14519_ (.A1(_06406_),
    .A2(_06513_),
    .B(_06514_),
    .ZN(_06515_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14520_ (.A1(_06479_),
    .A2(_06486_),
    .ZN(_06516_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _14521_ (.A1(_06476_),
    .A2(_06487_),
    .B(_06516_),
    .ZN(_06517_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _14522_ (.A1(_06412_),
    .A2(_06470_),
    .Z(_06518_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _14523_ (.A1(_06471_),
    .A2(_06488_),
    .B(_06518_),
    .ZN(_06519_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _14524_ (.I(_06484_),
    .Z(_06520_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _14525_ (.A1(_06520_),
    .A2(_06254_),
    .B(_06483_),
    .ZN(_06521_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14526_ (.A1(_06484_),
    .A2(_06254_),
    .A3(_06483_),
    .ZN(_06522_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _14527_ (.A1(_06480_),
    .A2(_06521_),
    .B(_06522_),
    .ZN(_06523_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14528_ (.A1(_06453_),
    .A2(_06467_),
    .ZN(_06524_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14529_ (.A1(_06450_),
    .A2(_06468_),
    .ZN(_06525_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14530_ (.A1(_06524_),
    .A2(_06525_),
    .ZN(_06526_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14531_ (.A1(_06484_),
    .A2(_04631_),
    .ZN(_06527_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _14532_ (.A1(_06455_),
    .A2(_06457_),
    .Z(_06528_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _14533_ (.A1(_06455_),
    .A2(_06457_),
    .Z(_06529_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _14534_ (.A1(_06454_),
    .A2(_06528_),
    .B(_06529_),
    .ZN(_06530_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14535_ (.A1(_06356_),
    .A2(_04667_),
    .ZN(_06531_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _14536_ (.A1(_06527_),
    .A2(_06530_),
    .A3(_06531_),
    .Z(_06532_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14537_ (.A1(_06526_),
    .A2(_06532_),
    .Z(_06533_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _14538_ (.A1(_06523_),
    .A2(_06533_),
    .ZN(_06534_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14539_ (.A1(_06415_),
    .A2(_06446_),
    .ZN(_06535_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14540_ (.A1(_06447_),
    .A2(_06469_),
    .ZN(_06536_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14541_ (.A1(_06535_),
    .A2(_06536_),
    .ZN(_06537_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14542_ (.A1(_06460_),
    .A2(_06465_),
    .ZN(_06538_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14543_ (.A1(_06458_),
    .A2(_06466_),
    .ZN(_06539_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14544_ (.A1(_06538_),
    .A2(_06539_),
    .ZN(_06540_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14545_ (.A1(_06438_),
    .A2(_06443_),
    .ZN(_06541_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _14546_ (.A1(_06435_),
    .A2(_06444_),
    .B(_06541_),
    .ZN(_06542_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14547_ (.A1(\filters.band[29] ),
    .A2(_05446_),
    .ZN(_06543_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14548_ (.A1(_06380_),
    .A2(_04600_),
    .ZN(_06544_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14549_ (.A1(\filters.band[30] ),
    .A2(_04506_),
    .ZN(_06545_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _14550_ (.A1(_06544_),
    .A2(_06545_),
    .Z(_06546_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14551_ (.A1(_06544_),
    .A2(_06545_),
    .ZN(_06547_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14552_ (.A1(_06546_),
    .A2(_06547_),
    .ZN(_06548_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14553_ (.A1(_06543_),
    .A2(_06548_),
    .Z(_06549_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14554_ (.A1(_06359_),
    .A2(_06093_),
    .A3(_06464_),
    .ZN(_06550_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _14555_ (.A1(_06462_),
    .A2(_06463_),
    .B(_06550_),
    .ZN(_06551_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14556_ (.A1(_04575_),
    .A2(_06008_),
    .ZN(_06552_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14557_ (.A1(_05512_),
    .A2(_05796_),
    .ZN(_06553_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14558_ (.A1(_05510_),
    .A2(_06005_),
    .ZN(_06554_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14559_ (.A1(_06553_),
    .A2(_06554_),
    .Z(_06555_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _14560_ (.A1(_06552_),
    .A2(_06555_),
    .ZN(_06556_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14561_ (.A1(_06551_),
    .A2(_06556_),
    .Z(_06557_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14562_ (.A1(_06549_),
    .A2(_06557_),
    .Z(_06558_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14563_ (.A1(_06542_),
    .A2(_06558_),
    .Z(_06559_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _14564_ (.A1(_06540_),
    .A2(_06559_),
    .ZN(_06560_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14565_ (.A1(_06417_),
    .A2(_06431_),
    .ZN(_06561_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14566_ (.A1(_06432_),
    .A2(_06445_),
    .ZN(_06562_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14567_ (.A1(_06561_),
    .A2(_06562_),
    .ZN(_06563_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14568_ (.A1(_04355_),
    .A2(_05775_),
    .A3(_06442_),
    .ZN(_06564_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _14569_ (.A1(_06440_),
    .A2(_06441_),
    .B(_06564_),
    .ZN(_06565_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14570_ (.A1(_04446_),
    .A2(_05449_),
    .A3(_06428_),
    .ZN(_06566_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _14571_ (.A1(_06426_),
    .A2(_06427_),
    .B(_06566_),
    .ZN(_06567_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14572_ (.A1(_04326_),
    .A2(_05891_),
    .ZN(_06568_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14573_ (.A1(_04452_),
    .A2(_05505_),
    .ZN(_06569_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14574_ (.A1(_04893_),
    .A2(_05687_),
    .ZN(_06570_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14575_ (.A1(_06569_),
    .A2(_06570_),
    .Z(_06571_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _14576_ (.A1(_06568_),
    .A2(_06571_),
    .ZN(_06572_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14577_ (.A1(_06567_),
    .A2(_06572_),
    .Z(_06573_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _14578_ (.A1(_06565_),
    .A2(_06573_),
    .ZN(_06574_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14579_ (.A1(_06420_),
    .A2(_06424_),
    .ZN(_06575_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _14580_ (.A1(_06425_),
    .A2(_06430_),
    .B(_06575_),
    .ZN(_06576_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14581_ (.A1(_04802_),
    .A2(_05501_),
    .ZN(_06577_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14582_ (.A1(_05909_),
    .A2(_05367_),
    .ZN(_06578_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14583_ (.A1(_04806_),
    .A2(_05448_),
    .ZN(_06579_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _14584_ (.A1(_06577_),
    .A2(_06578_),
    .A3(_06579_),
    .ZN(_06580_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _14585_ (.A1(_06421_),
    .A2(_06422_),
    .Z(_06581_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _14586_ (.A1(_06421_),
    .A2(_06422_),
    .Z(_06582_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _14587_ (.A1(_06581_),
    .A2(_06423_),
    .B(_06582_),
    .ZN(_06583_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14588_ (.A1(_04820_),
    .A2(_05280_),
    .ZN(_06584_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14589_ (.A1(_04924_),
    .A2(_05626_),
    .ZN(_06585_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14590_ (.A1(_05624_),
    .A2(_05091_),
    .ZN(_06586_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _14591_ (.A1(_06584_),
    .A2(_06585_),
    .A3(_06586_),
    .ZN(_06587_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14592_ (.A1(_06583_),
    .A2(_06587_),
    .Z(_06588_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _14593_ (.A1(_06576_),
    .A2(_06580_),
    .A3(_06588_),
    .Z(_06589_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _14594_ (.A1(_06574_),
    .A2(_06589_),
    .ZN(_06590_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _14595_ (.I(_06590_),
    .ZN(_06591_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14596_ (.A1(_06563_),
    .A2(_06591_),
    .Z(_06592_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _14597_ (.A1(_06560_),
    .A2(_06592_),
    .ZN(_06593_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14598_ (.A1(_06537_),
    .A2(_06593_),
    .Z(_06594_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _14599_ (.A1(_06534_),
    .A2(_06594_),
    .ZN(_06595_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _14600_ (.A1(_06519_),
    .A2(_06595_),
    .ZN(_06596_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _14601_ (.A1(_06517_),
    .A2(_06596_),
    .ZN(_06597_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14602_ (.A1(_06515_),
    .A2(_06597_),
    .Z(_06598_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _14603_ (.A1(_06512_),
    .A2(_06598_),
    .ZN(_06599_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14604_ (.A1(\filters.low[10] ),
    .A2(_03377_),
    .ZN(_06600_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _14605_ (.A1(_03396_),
    .A2(_06067_),
    .B(_06600_),
    .ZN(_06601_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _14606_ (.A1(_06599_),
    .A2(_06601_),
    .ZN(_06602_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _14607_ (.A1(_06400_),
    .A2(_06502_),
    .Z(_06603_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14608_ (.A1(_06499_),
    .A2(_06501_),
    .ZN(_06604_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14609_ (.A1(_06499_),
    .A2(_06501_),
    .ZN(_06605_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _14610_ (.A1(_06503_),
    .A2(_06604_),
    .B(_06605_),
    .ZN(_06606_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _14611_ (.A1(_06298_),
    .A2(_06603_),
    .B(_06606_),
    .ZN(_06607_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14612_ (.A1(_06602_),
    .A2(_06607_),
    .Z(_06608_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14613_ (.A1(_06403_),
    .A2(_06608_),
    .ZN(_06609_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _14614_ (.I(_06186_),
    .Z(_06610_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _14615_ (.A1(_03396_),
    .A2(_06508_),
    .B(_06609_),
    .C(_06610_),
    .ZN(_00536_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _14616_ (.I(_06519_),
    .ZN(_06611_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _14617_ (.A1(_06611_),
    .A2(_06595_),
    .Z(_06612_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _14618_ (.A1(_06517_),
    .A2(_06596_),
    .B(_06612_),
    .ZN(_06613_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _14619_ (.I(_06356_),
    .Z(_06614_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _14620_ (.A1(_06614_),
    .A2(_06473_),
    .B(_06530_),
    .ZN(_06615_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14621_ (.A1(_06356_),
    .A2(_06473_),
    .A3(_06530_),
    .ZN(_06616_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _14622_ (.A1(_06527_),
    .A2(_06615_),
    .B(_06616_),
    .ZN(_06617_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14623_ (.A1(_04222_),
    .A2(_06383_),
    .ZN(_06618_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14624_ (.A1(_06520_),
    .A2(_04601_),
    .ZN(_06619_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14625_ (.A1(_06567_),
    .A2(_06572_),
    .ZN(_06620_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14626_ (.A1(_06565_),
    .A2(_06573_),
    .ZN(_06621_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14627_ (.A1(_06620_),
    .A2(_06621_),
    .ZN(_06622_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14628_ (.A1(_05909_),
    .A2(_05561_),
    .ZN(_06623_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _14629_ (.A1(_06578_),
    .A2(_06579_),
    .Z(_06624_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _14630_ (.A1(_06578_),
    .A2(_06579_),
    .Z(_06625_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _14631_ (.A1(_06577_),
    .A2(_06624_),
    .B(_06625_),
    .ZN(_06626_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14632_ (.A1(_06623_),
    .A2(_06626_),
    .Z(_06627_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14633_ (.A1(_04318_),
    .A2(_05980_),
    .ZN(_06628_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14634_ (.A1(_04447_),
    .A2(_05766_),
    .ZN(_06629_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14635_ (.A1(_05624_),
    .A2(_05281_),
    .ZN(_06630_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _14636_ (.A1(_06585_),
    .A2(_06586_),
    .Z(_06631_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _14637_ (.A1(_06585_),
    .A2(_06586_),
    .Z(_06632_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _14638_ (.A1(_06584_),
    .A2(_06631_),
    .B(_06632_),
    .ZN(_06633_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _14639_ (.A1(_06629_),
    .A2(_06630_),
    .A3(_06633_),
    .Z(_06634_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _14640_ (.A1(_06627_),
    .A2(_06628_),
    .A3(_06634_),
    .Z(_06635_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _14641_ (.A1(_06619_),
    .A2(_06622_),
    .A3(_06635_),
    .Z(_06636_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _14642_ (.I(_06592_),
    .ZN(_06637_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14643_ (.A1(_06563_),
    .A2(_06591_),
    .ZN(_06638_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _14644_ (.A1(_06560_),
    .A2(_06637_),
    .B(_06638_),
    .ZN(_06639_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14645_ (.A1(_06472_),
    .A2(_04576_),
    .ZN(_06640_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14646_ (.A1(_04576_),
    .A2(_06383_),
    .A3(_06555_),
    .ZN(_06641_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _14647_ (.A1(_06553_),
    .A2(_06554_),
    .B(_06641_),
    .ZN(_06642_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14648_ (.A1(_05509_),
    .A2(_06096_),
    .ZN(_06643_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14649_ (.A1(_06551_),
    .A2(_06556_),
    .ZN(_06644_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14650_ (.A1(_06549_),
    .A2(_06557_),
    .ZN(_06645_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14651_ (.A1(_06644_),
    .A2(_06645_),
    .ZN(_06646_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14652_ (.A1(\filters.band[31] ),
    .A2(_04634_),
    .ZN(_06647_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _14653_ (.A1(_06643_),
    .A2(_06646_),
    .A3(_06647_),
    .Z(_06648_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _14654_ (.A1(_06640_),
    .A2(_06642_),
    .A3(_06648_),
    .Z(_06649_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14655_ (.A1(_06639_),
    .A2(_06649_),
    .Z(_06650_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _14656_ (.A1(_06618_),
    .A2(_06636_),
    .A3(_06650_),
    .Z(_06651_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _14657_ (.A1(_06613_),
    .A2(_06617_),
    .A3(_06651_),
    .Z(_06652_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14658_ (.A1(_06614_),
    .A2(_05982_),
    .ZN(_06653_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _14659_ (.A1(_06542_),
    .A2(_06558_),
    .Z(_06654_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _14660_ (.A1(_06540_),
    .A2(_06559_),
    .B(_06654_),
    .ZN(_06655_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14661_ (.A1(_06526_),
    .A2(_06532_),
    .ZN(_06656_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14662_ (.A1(_06523_),
    .A2(_06533_),
    .ZN(_06657_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14663_ (.A1(_06656_),
    .A2(_06657_),
    .ZN(_06658_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _14664_ (.I(_06594_),
    .ZN(_06659_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14665_ (.A1(_06537_),
    .A2(_06593_),
    .ZN(_06660_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _14666_ (.A1(_06534_),
    .A2(_06659_),
    .B(_06660_),
    .ZN(_06661_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _14667_ (.A1(_06655_),
    .A2(_06658_),
    .A3(_06661_),
    .Z(_06662_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14668_ (.A1(_06456_),
    .A2(_06473_),
    .ZN(_06663_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14669_ (.A1(_06332_),
    .A2(_06086_),
    .ZN(_06664_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _14670_ (.A1(_06580_),
    .A2(_06588_),
    .Z(_06665_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14671_ (.A1(_06580_),
    .A2(_06588_),
    .ZN(_06666_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _14672_ (.A1(_06576_),
    .A2(_06665_),
    .A3(_06666_),
    .B1(_06589_),
    .B2(_06574_),
    .ZN(_06667_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14673_ (.A1(_04806_),
    .A2(_05663_),
    .ZN(_06668_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14674_ (.A1(_04820_),
    .A2(_05370_),
    .ZN(_06669_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14675_ (.A1(_05268_),
    .A2(_05626_),
    .ZN(_06670_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14676_ (.A1(_06583_),
    .A2(_06587_),
    .ZN(_06671_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14677_ (.A1(_06580_),
    .A2(_06588_),
    .ZN(_06672_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14678_ (.A1(_06671_),
    .A2(_06672_),
    .ZN(_06673_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _14679_ (.A1(_06669_),
    .A2(_06670_),
    .A3(_06673_),
    .Z(_06674_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14680_ (.A1(\filters.band[30] ),
    .A2(_04633_),
    .ZN(_06675_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14681_ (.A1(_06332_),
    .A2(_05980_),
    .A3(_06571_),
    .ZN(_06676_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _14682_ (.A1(_04453_),
    .A2(_05883_),
    .Z(_06677_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14683_ (.A1(_06441_),
    .A2(_06676_),
    .A3(_06677_),
    .ZN(_06678_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _14684_ (.A1(_06676_),
    .A2(_06677_),
    .B(_06678_),
    .ZN(_06679_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14685_ (.A1(_06675_),
    .A2(_06679_),
    .Z(_06680_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _14686_ (.A1(_06668_),
    .A2(_06674_),
    .A3(_06680_),
    .Z(_06681_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _14687_ (.A1(_06664_),
    .A2(_06667_),
    .A3(_06681_),
    .Z(_06682_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _14688_ (.A1(_06543_),
    .A2(_06548_),
    .B(_06546_),
    .ZN(_06683_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _14689_ (.A1(_06663_),
    .A2(_06682_),
    .A3(_06683_),
    .Z(_06684_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _14690_ (.A1(_06653_),
    .A2(_06662_),
    .A3(_06684_),
    .Z(_06685_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14691_ (.A1(_06515_),
    .A2(_06597_),
    .ZN(_06686_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _14692_ (.A1(_06512_),
    .A2(_06598_),
    .B(_06686_),
    .ZN(_06687_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _14693_ (.A1(_06652_),
    .A2(_06685_),
    .A3(_06687_),
    .Z(_06688_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _14694_ (.I(_06688_),
    .Z(_06689_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14695_ (.A1(_03411_),
    .A2(_03221_),
    .ZN(_06690_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _14696_ (.A1(_03412_),
    .A2(_03378_),
    .B(_06690_),
    .ZN(_06691_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _14697_ (.A1(_06689_),
    .A2(_06691_),
    .ZN(_06692_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14698_ (.A1(_06599_),
    .A2(_06601_),
    .ZN(_06693_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _14699_ (.A1(_06602_),
    .A2(_06607_),
    .B(_06693_),
    .ZN(_06694_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14700_ (.A1(_06692_),
    .A2(_06694_),
    .Z(_06695_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _14701_ (.A1(\filters.band[11] ),
    .A2(_05540_),
    .B(_05541_),
    .ZN(_06696_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _14702_ (.A1(_04161_),
    .A2(_06695_),
    .B(_06696_),
    .ZN(_00537_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14703_ (.A1(_06400_),
    .A2(_06502_),
    .ZN(_06697_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _14704_ (.A1(_06602_),
    .A2(_06697_),
    .A3(_06692_),
    .ZN(_06698_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _14705_ (.I(_06602_),
    .ZN(_06699_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _14706_ (.I(_06688_),
    .Z(_06700_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _14707_ (.I(_06700_),
    .Z(_06701_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _14708_ (.A1(_06701_),
    .A2(_06691_),
    .ZN(_06702_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _14709_ (.I(_06700_),
    .Z(_06703_));
 gf180mcu_fd_sc_mcu7t5v0__or2_4 _14710_ (.A1(_06703_),
    .A2(_06691_),
    .Z(_06704_));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 _14711_ (.A1(_06699_),
    .A2(_06606_),
    .A3(_06702_),
    .A4(_06704_),
    .Z(_06705_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _14712_ (.I(_06700_),
    .Z(_06706_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _14713_ (.A1(_06706_),
    .A2(_06691_),
    .ZN(_06707_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _14714_ (.A1(_06693_),
    .A2(_06707_),
    .B(_06702_),
    .ZN(_06708_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _14715_ (.A1(_06298_),
    .A2(_06698_),
    .B(_06705_),
    .C(_06708_),
    .ZN(_06709_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _14716_ (.I(_06067_),
    .Z(_06710_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14717_ (.A1(_03422_),
    .A2(_06397_),
    .ZN(_06711_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _14718_ (.A1(_03423_),
    .A2(_06710_),
    .B(_06711_),
    .ZN(_06712_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14719_ (.A1(_06689_),
    .A2(_06712_),
    .Z(_06713_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14720_ (.A1(net30),
    .A2(_06713_),
    .Z(_06714_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _14721_ (.A1(\filters.band[12] ),
    .A2(_05540_),
    .B(_05541_),
    .ZN(_06715_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _14722_ (.A1(_04161_),
    .A2(_06714_),
    .B(_06715_),
    .ZN(_00538_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _14723_ (.I(_06703_),
    .Z(_06716_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _14724_ (.I(_06716_),
    .Z(_06717_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _14725_ (.I(_06717_),
    .Z(_06718_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14726_ (.I(_06718_),
    .Z(_06719_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _14727_ (.I(_06719_),
    .Z(_06720_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14728_ (.A1(_06720_),
    .A2(_06712_),
    .ZN(_06721_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _14729_ (.I(_06719_),
    .Z(_06722_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14730_ (.A1(_06722_),
    .A2(_06712_),
    .ZN(_06723_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _14731_ (.A1(net30),
    .A2(_06721_),
    .B(_06723_),
    .ZN(_06724_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14732_ (.A1(_03439_),
    .A2(_06710_),
    .ZN(_06725_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _14733_ (.A1(_03440_),
    .A2(_03222_),
    .B(_06725_),
    .ZN(_06726_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14734_ (.A1(_06689_),
    .A2(_06726_),
    .Z(_06727_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14735_ (.A1(_06724_),
    .A2(_06727_),
    .Z(_06728_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14736_ (.A1(_06403_),
    .A2(_06728_),
    .ZN(_06729_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _14737_ (.A1(_03440_),
    .A2(_06508_),
    .B(_06729_),
    .C(_06610_),
    .ZN(_00539_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14738_ (.A1(_03455_),
    .A2(_06397_),
    .ZN(_06730_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _14739_ (.A1(_03456_),
    .A2(_03222_),
    .B(_06730_),
    .ZN(_06731_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _14740_ (.A1(_06703_),
    .A2(_06731_),
    .Z(_06732_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14741_ (.A1(_06713_),
    .A2(_06727_),
    .ZN(_06733_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _14742_ (.I(_06716_),
    .Z(_06734_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _14743_ (.A1(_06712_),
    .A2(_06726_),
    .B(_06734_),
    .ZN(_06735_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _14744_ (.A1(net30),
    .A2(_06733_),
    .B(_06735_),
    .ZN(_06736_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14745_ (.A1(_06732_),
    .A2(_06736_),
    .Z(_06737_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14746_ (.A1(_06403_),
    .A2(_06737_),
    .ZN(_06738_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _14747_ (.A1(_03456_),
    .A2(_06508_),
    .B(_06738_),
    .C(_06610_),
    .ZN(_00540_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _14748_ (.I(\filters.band[15] ),
    .ZN(_06739_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14749_ (.A1(_03468_),
    .A2(_06710_),
    .ZN(_06740_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _14750_ (.A1(_06739_),
    .A2(_03222_),
    .B(_06740_),
    .ZN(_06741_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14751_ (.A1(_06741_),
    .A2(_06703_),
    .Z(_06742_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14752_ (.A1(_06722_),
    .A2(_06731_),
    .ZN(_06743_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14753_ (.A1(_06732_),
    .A2(_06736_),
    .ZN(_06744_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14754_ (.A1(_06743_),
    .A2(_06744_),
    .ZN(_06745_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14755_ (.A1(_06742_),
    .A2(_06745_),
    .Z(_06746_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14756_ (.A1(_05544_),
    .A2(_06746_),
    .ZN(_06747_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _14757_ (.A1(_06739_),
    .A2(_06508_),
    .B(_06747_),
    .C(_06610_),
    .ZN(_00541_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14758_ (.I(_05546_),
    .Z(_06748_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _14759_ (.A1(_06732_),
    .A2(_06742_),
    .ZN(_06749_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _14760_ (.A1(_06749_),
    .A2(_06733_),
    .Z(_06750_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _14761_ (.A1(_06731_),
    .A2(_06741_),
    .B(_06734_),
    .ZN(_06751_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _14762_ (.A1(_06735_),
    .A2(_06749_),
    .B1(_06750_),
    .B2(_06709_),
    .C(_06751_),
    .ZN(_06752_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _14763_ (.I(_06752_),
    .Z(_06753_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _14764_ (.I(_06700_),
    .Z(_06754_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _14765_ (.I(_03472_),
    .Z(_06755_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _14766_ (.I0(\filters.low[16] ),
    .I1(\filters.band[16] ),
    .S(_06755_),
    .Z(_06756_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _14767_ (.A1(_06754_),
    .A2(_06756_),
    .Z(_06757_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14768_ (.A1(_06753_),
    .A2(_06757_),
    .Z(_06758_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14769_ (.A1(_06748_),
    .A2(_06758_),
    .ZN(_06759_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14770_ (.I(_04159_),
    .Z(_06760_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _14771_ (.I(_06760_),
    .Z(_06761_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _14772_ (.I(_03733_),
    .Z(_06762_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14773_ (.I(_06762_),
    .Z(_06763_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _14774_ (.A1(\filters.band[16] ),
    .A2(_06761_),
    .B(_06763_),
    .ZN(_06764_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14775_ (.A1(_06759_),
    .A2(_06764_),
    .ZN(_00542_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _14776_ (.I(_06716_),
    .Z(_06765_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _14777_ (.I(_06765_),
    .Z(_06766_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14778_ (.I(_06766_),
    .Z(_06767_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _14779_ (.I(_06767_),
    .Z(_06768_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _14780_ (.I(_06768_),
    .Z(_06769_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _14781_ (.A1(_06769_),
    .A2(_06756_),
    .Z(_06770_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _14782_ (.A1(_06753_),
    .A2(_06757_),
    .B(_06770_),
    .ZN(_06771_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _14783_ (.I0(\filters.low[17] ),
    .I1(\filters.band[17] ),
    .S(_06755_),
    .Z(_06772_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14784_ (.A1(_06754_),
    .A2(_06772_),
    .Z(_06773_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14785_ (.A1(_06771_),
    .A2(_06773_),
    .Z(_06774_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _14786_ (.I(_03721_),
    .Z(_06775_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _14787_ (.A1(\filters.band[17] ),
    .A2(_04160_),
    .B(_06775_),
    .ZN(_06776_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _14788_ (.A1(_06761_),
    .A2(_06774_),
    .B(_06776_),
    .ZN(_00543_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _14789_ (.I(_06689_),
    .Z(_06777_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _14790_ (.I0(\filters.low[18] ),
    .I1(\filters.band[18] ),
    .S(_06073_),
    .Z(_06778_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _14791_ (.A1(_06777_),
    .A2(_06778_),
    .ZN(_06779_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _14792_ (.A1(_06756_),
    .A2(_06772_),
    .B(_06765_),
    .ZN(_06780_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14793_ (.A1(_06753_),
    .A2(_06757_),
    .A3(_06773_),
    .ZN(_06781_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14794_ (.A1(_06780_),
    .A2(_06781_),
    .ZN(_06782_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _14795_ (.A1(_06779_),
    .A2(_06782_),
    .ZN(_06783_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14796_ (.A1(_06748_),
    .A2(_06783_),
    .ZN(_06784_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14797_ (.I(_06760_),
    .Z(_06785_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _14798_ (.A1(\filters.band[18] ),
    .A2(_06785_),
    .B(_06763_),
    .ZN(_06786_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14799_ (.A1(_06784_),
    .A2(_06786_),
    .ZN(_00544_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _14800_ (.I0(\filters.low[19] ),
    .I1(\filters.band[19] ),
    .S(_06755_),
    .Z(_06787_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _14801_ (.A1(_06706_),
    .A2(_06787_),
    .ZN(_06788_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _14802_ (.A1(_06780_),
    .A2(_06781_),
    .B(_06779_),
    .ZN(_06789_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _14803_ (.A1(_06769_),
    .A2(_06778_),
    .B(_06789_),
    .ZN(_06790_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14804_ (.A1(_06788_),
    .A2(_06790_),
    .Z(_06791_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14805_ (.A1(_06748_),
    .A2(_06791_),
    .ZN(_06792_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _14806_ (.A1(\filters.band[19] ),
    .A2(_06785_),
    .B(_06763_),
    .ZN(_06793_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14807_ (.A1(_06792_),
    .A2(_06793_),
    .ZN(_00545_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _14808_ (.I0(\filters.low[20] ),
    .I1(\filters.band[20] ),
    .S(_03472_),
    .Z(_06794_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _14809_ (.A1(_06701_),
    .A2(_06794_),
    .ZN(_06795_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14810_ (.A1(_06757_),
    .A2(_06773_),
    .ZN(_06796_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _14811_ (.A1(_06779_),
    .A2(_06796_),
    .A3(_06788_),
    .ZN(_06797_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _14812_ (.A1(_06778_),
    .A2(_06787_),
    .B(_06734_),
    .ZN(_06798_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_4 _14813_ (.A1(_06779_),
    .A2(_06780_),
    .A3(_06788_),
    .B(_06798_),
    .ZN(_06799_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _14814_ (.A1(_06753_),
    .A2(_06797_),
    .B(_06799_),
    .ZN(_06800_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14815_ (.A1(_06795_),
    .A2(_06800_),
    .Z(_06801_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14816_ (.A1(_06748_),
    .A2(_06801_),
    .ZN(_06802_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _14817_ (.A1(\filters.band[20] ),
    .A2(_06785_),
    .B(_06763_),
    .ZN(_06803_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14818_ (.A1(_06802_),
    .A2(_06803_),
    .ZN(_00546_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14819_ (.I(_05546_),
    .Z(_06804_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14820_ (.A1(_06795_),
    .A2(_06800_),
    .ZN(_06805_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _14821_ (.A1(_06769_),
    .A2(_06794_),
    .B(_06805_),
    .ZN(_06806_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _14822_ (.I0(\filters.low[21] ),
    .I1(\filters.band[21] ),
    .S(_06073_),
    .Z(_06807_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _14823_ (.A1(_06777_),
    .A2(_06807_),
    .ZN(_06808_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14824_ (.A1(_06806_),
    .A2(_06808_),
    .Z(_06809_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14825_ (.A1(_06804_),
    .A2(_06809_),
    .ZN(_06810_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14826_ (.I(_06762_),
    .Z(_06811_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _14827_ (.A1(\filters.band[21] ),
    .A2(_06785_),
    .B(_06811_),
    .ZN(_06812_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14828_ (.A1(_06810_),
    .A2(_06812_),
    .ZN(_00547_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _14829_ (.I0(\filters.low[22] ),
    .I1(\filters.band[22] ),
    .S(_06073_),
    .Z(_06813_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _14830_ (.A1(_06777_),
    .A2(_06813_),
    .ZN(_06814_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _14831_ (.I(_06814_),
    .ZN(_06815_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _14832_ (.A1(_06794_),
    .A2(_06807_),
    .B(_06765_),
    .ZN(_06816_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _14833_ (.A1(_06795_),
    .A2(_06800_),
    .A3(_06808_),
    .B(_06816_),
    .ZN(_06817_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14834_ (.A1(_06815_),
    .A2(_06817_),
    .Z(_06818_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14835_ (.A1(_06804_),
    .A2(_06818_),
    .ZN(_06819_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14836_ (.I(_06760_),
    .Z(_06820_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _14837_ (.A1(\filters.band[22] ),
    .A2(_06820_),
    .B(_06811_),
    .ZN(_06821_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14838_ (.A1(_06819_),
    .A2(_06821_),
    .ZN(_00548_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _14839_ (.I(\filters.low[23] ),
    .ZN(_06822_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14840_ (.A1(\filters.band[23] ),
    .A2(_06755_),
    .ZN(_06823_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _14841_ (.A1(_06822_),
    .A2(_03473_),
    .B(_06823_),
    .ZN(_06824_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _14842_ (.A1(_06777_),
    .A2(_06824_),
    .ZN(_06825_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _14843_ (.A1(_06720_),
    .A2(_06813_),
    .Z(_06826_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _14844_ (.A1(_06815_),
    .A2(_06817_),
    .B(_06826_),
    .ZN(_06827_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14845_ (.A1(_06825_),
    .A2(_06827_),
    .Z(_06828_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14846_ (.A1(_06804_),
    .A2(_06828_),
    .ZN(_06829_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _14847_ (.A1(\filters.band[23] ),
    .A2(_06820_),
    .B(_06811_),
    .ZN(_06830_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14848_ (.A1(_06829_),
    .A2(_06830_),
    .ZN(_00549_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _14849_ (.A1(_06795_),
    .A2(_06808_),
    .A3(_06814_),
    .A4(_06825_),
    .ZN(_06831_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _14850_ (.A1(_06797_),
    .A2(_06831_),
    .Z(_06832_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _14851_ (.A1(_06813_),
    .A2(_06824_),
    .B(_06717_),
    .ZN(_06833_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _14852_ (.A1(_06814_),
    .A2(_06816_),
    .A3(_06825_),
    .B(_06833_),
    .ZN(_06834_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _14853_ (.A1(_06799_),
    .A2(_06831_),
    .B1(_06832_),
    .B2(_06752_),
    .C(_06834_),
    .ZN(_06835_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _14854_ (.I(_06701_),
    .Z(_06836_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _14855_ (.I(\filters.low[24] ),
    .ZN(_06837_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14856_ (.A1(\filters.band[24] ),
    .A2(_03474_),
    .ZN(_06838_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _14857_ (.A1(_06837_),
    .A2(_03474_),
    .B(_06838_),
    .ZN(_06839_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14858_ (.A1(_06836_),
    .A2(_06839_),
    .Z(_06840_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14859_ (.A1(_06835_),
    .A2(_06840_),
    .Z(_06841_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _14860_ (.A1(\filters.band[24] ),
    .A2(_04160_),
    .B(_06775_),
    .ZN(_06842_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _14861_ (.A1(_06761_),
    .A2(_06841_),
    .B(_06842_),
    .ZN(_00550_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _14862_ (.I(_06840_),
    .ZN(_06843_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14863_ (.A1(_06722_),
    .A2(_06839_),
    .ZN(_06844_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _14864_ (.A1(_06835_),
    .A2(_06843_),
    .B(_06844_),
    .ZN(_06845_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _14865_ (.I0(\filters.low[25] ),
    .I1(\filters.band[25] ),
    .S(_03473_),
    .Z(_06846_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14866_ (.A1(_06836_),
    .A2(_06846_),
    .Z(_06847_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14867_ (.A1(_06845_),
    .A2(_06847_),
    .Z(_06848_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14868_ (.A1(_06804_),
    .A2(_06848_),
    .ZN(_06849_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _14869_ (.A1(\filters.band[25] ),
    .A2(_06820_),
    .B(_06811_),
    .ZN(_06850_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14870_ (.A1(_06849_),
    .A2(_06850_),
    .ZN(_00551_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14871_ (.I(_05546_),
    .Z(_06851_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _14872_ (.I(_06706_),
    .Z(_06852_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _14873_ (.I0(\filters.low[26] ),
    .I1(_06472_),
    .S(_03473_),
    .Z(_06853_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14874_ (.A1(_06852_),
    .A2(_06853_),
    .Z(_06854_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14875_ (.A1(_06840_),
    .A2(_06847_),
    .ZN(_06855_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _14876_ (.A1(_06839_),
    .A2(_06846_),
    .B(_06718_),
    .ZN(_06856_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _14877_ (.A1(net32),
    .A2(_06855_),
    .B(_06856_),
    .ZN(_06857_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14878_ (.A1(_06854_),
    .A2(_06857_),
    .Z(_06858_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14879_ (.A1(_06851_),
    .A2(_06858_),
    .ZN(_06859_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14880_ (.I(_06762_),
    .Z(_06860_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _14881_ (.A1(_06472_),
    .A2(_06820_),
    .B(_06860_),
    .ZN(_06861_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14882_ (.A1(_06859_),
    .A2(_06861_),
    .ZN(_00552_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _14883_ (.I(_06706_),
    .Z(_06862_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _14884_ (.I0(\filters.low[27] ),
    .I1(_06520_),
    .S(_03474_),
    .Z(_06863_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14885_ (.A1(_06862_),
    .A2(_06863_),
    .Z(_06864_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _14886_ (.A1(_06768_),
    .A2(_06853_),
    .Z(_06865_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _14887_ (.A1(_06854_),
    .A2(_06857_),
    .B(_06865_),
    .ZN(_06866_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _14888_ (.A1(_06864_),
    .A2(_06866_),
    .ZN(_06867_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14889_ (.A1(_06851_),
    .A2(_06867_),
    .ZN(_06868_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14890_ (.I(_06760_),
    .Z(_06869_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _14891_ (.A1(_06520_),
    .A2(_06869_),
    .B(_06860_),
    .ZN(_06870_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14892_ (.A1(_06868_),
    .A2(_06870_),
    .ZN(_00553_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _14893_ (.A1(_06854_),
    .A2(_06864_),
    .ZN(_06871_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _14894_ (.A1(_06855_),
    .A2(_06871_),
    .Z(_06872_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _14895_ (.A1(_06853_),
    .A2(_06863_),
    .B(_06718_),
    .ZN(_06873_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _14896_ (.A1(_06856_),
    .A2(_06871_),
    .B1(_06872_),
    .B2(_06835_),
    .C(_06873_),
    .ZN(_06874_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _14897_ (.I(\filters.low[28] ),
    .ZN(_06875_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14898_ (.A1(_06614_),
    .A2(_03475_),
    .ZN(_06876_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _14899_ (.A1(_06875_),
    .A2(_03476_),
    .B(_06876_),
    .ZN(_06877_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14900_ (.A1(_06766_),
    .A2(_06877_),
    .Z(_06878_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14901_ (.A1(_06874_),
    .A2(_06878_),
    .Z(_06879_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14902_ (.A1(_06851_),
    .A2(_06879_),
    .ZN(_06880_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _14903_ (.A1(_06614_),
    .A2(_06869_),
    .B(_06860_),
    .ZN(_06881_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14904_ (.A1(_06880_),
    .A2(_06881_),
    .ZN(_00554_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _14905_ (.I(\filters.low[29] ),
    .ZN(_06882_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14906_ (.A1(_06456_),
    .A2(_03475_),
    .ZN(_06883_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _14907_ (.A1(_06882_),
    .A2(_03475_),
    .B(_06883_),
    .ZN(_06884_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _14908_ (.A1(_06718_),
    .A2(_06884_),
    .ZN(_06885_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _14909_ (.A1(_06719_),
    .A2(_06877_),
    .Z(_06886_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _14910_ (.A1(_06874_),
    .A2(_06878_),
    .B(_06886_),
    .ZN(_06887_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14911_ (.A1(_06885_),
    .A2(_06887_),
    .Z(_06888_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14912_ (.A1(_06851_),
    .A2(_06888_),
    .ZN(_06889_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _14913_ (.A1(_06456_),
    .A2(_06869_),
    .B(_06860_),
    .ZN(_06890_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14914_ (.A1(_06889_),
    .A2(_06890_),
    .ZN(_00555_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _14915_ (.I(\filters.low[30] ),
    .ZN(_06891_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14916_ (.A1(\filters.band[30] ),
    .A2(_03476_),
    .ZN(_06892_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _14917_ (.A1(_06891_),
    .A2(_03477_),
    .B(_06892_),
    .ZN(_06893_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _14918_ (.I(_06878_),
    .ZN(_06894_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _14919_ (.A1(_06894_),
    .A2(_06885_),
    .ZN(_06895_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _14920_ (.A1(_06768_),
    .A2(_06884_),
    .B1(_06895_),
    .B2(_06874_),
    .C(_06886_),
    .ZN(_06896_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _14921_ (.A1(_06722_),
    .A2(_06893_),
    .A3(net70),
    .ZN(_06897_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14922_ (.A1(_05547_),
    .A2(_06897_),
    .ZN(_06898_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _14923_ (.I(_06762_),
    .Z(_06899_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _14924_ (.A1(\filters.band[30] ),
    .A2(_06869_),
    .B(_06899_),
    .ZN(_06900_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14925_ (.A1(_06898_),
    .A2(_06900_),
    .ZN(_00556_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14926_ (.A1(_06720_),
    .A2(_06893_),
    .ZN(_06901_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14927_ (.A1(_06720_),
    .A2(_06893_),
    .ZN(_06902_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _14928_ (.A1(_06901_),
    .A2(_06896_),
    .B(_06902_),
    .ZN(_06903_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _14929_ (.I0(\filters.low[31] ),
    .I1(\filters.band[31] ),
    .S(_03477_),
    .Z(_06904_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _14930_ (.A1(_06769_),
    .A2(_06903_),
    .A3(_06904_),
    .ZN(_06905_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _14931_ (.A1(\filters.band[31] ),
    .A2(_04160_),
    .B(_06775_),
    .ZN(_06906_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _14932_ (.A1(_06761_),
    .A2(_06905_),
    .B(_06906_),
    .ZN(_00557_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14933_ (.A1(_03730_),
    .A2(_04170_),
    .ZN(_06907_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _14934_ (.I(_06907_),
    .Z(_06908_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _14935_ (.I(_06908_),
    .Z(_06909_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _14936_ (.I(_06909_),
    .Z(_06910_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _14937_ (.I(\filters.low[0] ),
    .ZN(_06911_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14938_ (.A1(_04558_),
    .A2(_04690_),
    .Z(_06912_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _14939_ (.I(_06908_),
    .Z(_06913_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _14940_ (.A1(_06911_),
    .A2(_06912_),
    .B(_06913_),
    .ZN(_06914_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _14941_ (.A1(_04558_),
    .A2(_04690_),
    .ZN(_06915_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14942_ (.A1(_05534_),
    .A2(_06915_),
    .ZN(_06916_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _14943_ (.I(_02353_),
    .Z(_06917_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _14944_ (.A1(_04214_),
    .A2(_06910_),
    .B1(_06914_),
    .B2(_06916_),
    .C(_06917_),
    .ZN(_00558_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14945_ (.I(_01932_),
    .Z(_06918_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _14946_ (.I(_06908_),
    .Z(_06919_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _14947_ (.A1(_04558_),
    .A2(_04690_),
    .B(_04691_),
    .ZN(_06920_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _14948_ (.A1(_04431_),
    .A2(_04519_),
    .A3(_06920_),
    .ZN(_06921_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _14949_ (.A1(_01759_),
    .A2(_01745_),
    .A3(\channels.sample1[0] ),
    .A4(\channels.sample2[0] ),
    .Z(_06922_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _14950_ (.A1(_01745_),
    .A2(\channels.sample1[0] ),
    .B1(\channels.sample2[0] ),
    .B2(_01759_),
    .ZN(_06923_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14951_ (.A1(_06922_),
    .A2(_06923_),
    .ZN(_06924_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14952_ (.A1(_01768_),
    .A2(\channels.sample3[0] ),
    .ZN(_06925_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _14953_ (.A1(_05647_),
    .A2(_06924_),
    .A3(_06925_),
    .ZN(_06926_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _14954_ (.I(_06926_),
    .ZN(_06927_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _14955_ (.A1(_06911_),
    .A2(_06912_),
    .B(_06927_),
    .ZN(_06928_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14956_ (.A1(_05534_),
    .A2(_06915_),
    .A3(_06926_),
    .ZN(_06929_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14957_ (.A1(_06921_),
    .A2(_06928_),
    .A3(_06929_),
    .ZN(_06930_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _14958_ (.A1(_06928_),
    .A2(_06929_),
    .B(_06921_),
    .ZN(_06931_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14959_ (.A1(_06909_),
    .A2(_06931_),
    .ZN(_06932_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _14960_ (.A1(\filters.high[1] ),
    .A2(_06919_),
    .B1(_06930_),
    .B2(_06932_),
    .ZN(_06933_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14961_ (.A1(_06918_),
    .A2(_06933_),
    .ZN(_00559_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _14962_ (.I(_06908_),
    .Z(_06934_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _14963_ (.A1(_06928_),
    .A2(_06930_),
    .Z(_06935_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _14964_ (.A1(_06922_),
    .A2(_06923_),
    .B(_06925_),
    .ZN(_06936_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14965_ (.A1(_01773_),
    .A2(\channels.sample3[0] ),
    .A3(_06924_),
    .ZN(_06937_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _14966_ (.A1(_05647_),
    .A2(_06936_),
    .A3(_06937_),
    .ZN(_06938_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _14967_ (.A1(_04520_),
    .A2(_04692_),
    .ZN(_06939_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _14968_ (.A1(_01758_),
    .A2(_01744_),
    .A3(\channels.sample1[1] ),
    .A4(\channels.sample2[1] ),
    .Z(_06940_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _14969_ (.A1(_01744_),
    .A2(\channels.sample1[1] ),
    .B1(\channels.sample2[1] ),
    .B2(_01758_),
    .ZN(_06941_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14970_ (.A1(_06940_),
    .A2(_06941_),
    .ZN(_06942_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14971_ (.A1(_01768_),
    .A2(\channels.sample3[1] ),
    .ZN(_06943_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14972_ (.A1(_06942_),
    .A2(_06943_),
    .Z(_06944_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _14973_ (.A1(_06922_),
    .A2(_06923_),
    .A3(_06925_),
    .ZN(_06945_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _14974_ (.A1(_06922_),
    .A2(_06945_),
    .ZN(_06946_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14975_ (.A1(_06944_),
    .A2(_06946_),
    .Z(_06947_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14976_ (.A1(\filters.low[2] ),
    .A2(_06947_),
    .Z(_06948_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _14977_ (.A1(_06939_),
    .A2(_05035_),
    .A3(_06948_),
    .Z(_06949_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _14978_ (.A1(_06938_),
    .A2(_06949_),
    .ZN(_06950_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _14979_ (.A1(_06935_),
    .A2(_06950_),
    .Z(_06951_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _14980_ (.I(_06907_),
    .Z(_06952_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _14981_ (.A1(_06935_),
    .A2(_06950_),
    .B(_06952_),
    .ZN(_06953_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _14982_ (.A1(\filters.high[2] ),
    .A2(_06934_),
    .B1(_06951_),
    .B2(_06953_),
    .ZN(_06954_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14983_ (.A1(_06918_),
    .A2(_06954_),
    .ZN(_00560_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _14984_ (.I(_06952_),
    .Z(_06955_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14985_ (.A1(\filters.high[3] ),
    .A2(_06955_),
    .ZN(_06956_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14986_ (.A1(_06938_),
    .A2(_06949_),
    .ZN(_06957_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _14987_ (.A1(_06935_),
    .A2(_06950_),
    .B(_06957_),
    .ZN(_06958_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14988_ (.A1(_06944_),
    .A2(_06946_),
    .ZN(_06959_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _14989_ (.I(_06943_),
    .ZN(_06960_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _14990_ (.A1(_06942_),
    .A2(_06960_),
    .B(_06940_),
    .ZN(_06961_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _14991_ (.A1(\filters.filt_2 ),
    .A2(\filters.filt_1 ),
    .A3(\channels.sample1[2] ),
    .A4(\channels.sample2[2] ),
    .Z(_06962_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _14992_ (.A1(\filters.filt_1 ),
    .A2(\channels.sample1[2] ),
    .B1(\channels.sample2[2] ),
    .B2(\filters.filt_2 ),
    .ZN(_06963_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _14993_ (.A1(_06962_),
    .A2(_06963_),
    .Z(_06964_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14994_ (.A1(\filters.filt_3 ),
    .A2(\channels.sample3[2] ),
    .ZN(_06965_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _14995_ (.A1(_06964_),
    .A2(_06965_),
    .ZN(_06966_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _14996_ (.A1(_06961_),
    .A2(_06966_),
    .ZN(_06967_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _14997_ (.A1(_06959_),
    .A2(_06967_),
    .ZN(_06968_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14998_ (.A1(\filters.low[3] ),
    .A2(_06968_),
    .Z(_06969_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _14999_ (.A1(_06939_),
    .A2(_05035_),
    .B(_05040_),
    .ZN(_06970_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _15000_ (.A1(net37),
    .A2(_06969_),
    .A3(_06970_),
    .Z(_06971_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _15001_ (.A1(_06939_),
    .A2(_05035_),
    .Z(_06972_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15002_ (.A1(_03268_),
    .A2(_06947_),
    .ZN(_06973_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15003_ (.A1(_06948_),
    .A2(_06972_),
    .B(_06973_),
    .ZN(_06974_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _15004_ (.A1(_06971_),
    .A2(_06974_),
    .Z(_06975_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15005_ (.A1(_06958_),
    .A2(_06975_),
    .B(_06952_),
    .ZN(_06976_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15006_ (.A1(_06958_),
    .A2(_06975_),
    .B(_06976_),
    .ZN(_06977_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15007_ (.I(_03940_),
    .Z(_06978_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _15008_ (.I(_06978_),
    .Z(_06979_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15009_ (.A1(_06956_),
    .A2(_06977_),
    .B(_06979_),
    .ZN(_00561_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15010_ (.A1(\filters.high[4] ),
    .A2(_06955_),
    .ZN(_06980_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15011_ (.A1(_04158_),
    .A2(_04776_),
    .ZN(_06981_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15012_ (.I(_06981_),
    .Z(_06982_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _15013_ (.I(_06982_),
    .Z(_06983_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _15014_ (.A1(_06944_),
    .A2(_06946_),
    .A3(_06967_),
    .B1(_06966_),
    .B2(_06961_),
    .ZN(_06984_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15015_ (.A1(_06964_),
    .A2(_06965_),
    .ZN(_06985_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15016_ (.A1(_06962_),
    .A2(_06985_),
    .ZN(_06986_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _15017_ (.A1(\filters.filt_2 ),
    .A2(\filters.filt_1 ),
    .A3(\channels.sample1[3] ),
    .A4(\channels.sample2[3] ),
    .Z(_06987_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _15018_ (.A1(_01744_),
    .A2(\channels.sample1[3] ),
    .B1(\channels.sample2[3] ),
    .B2(_01758_),
    .ZN(_06988_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _15019_ (.A1(_06987_),
    .A2(_06988_),
    .Z(_06989_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15020_ (.A1(_01768_),
    .A2(\channels.sample3[3] ),
    .ZN(_06990_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _15021_ (.A1(_06989_),
    .A2(_06990_),
    .ZN(_06991_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _15022_ (.A1(_06986_),
    .A2(_06991_),
    .Z(_06992_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _15023_ (.A1(_06984_),
    .A2(_06992_),
    .Z(_06993_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _15024_ (.I(_05016_),
    .ZN(_06994_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _15025_ (.A1(_04693_),
    .A2(_05036_),
    .B(_05042_),
    .ZN(_06995_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _15026_ (.A1(_06994_),
    .A2(_06995_),
    .Z(_06996_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _15027_ (.A1(\filters.low[4] ),
    .A2(_06993_),
    .A3(_06996_),
    .ZN(_06997_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _15028_ (.A1(net38),
    .A2(_06970_),
    .ZN(_06998_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15029_ (.A1(_03282_),
    .A2(_06968_),
    .ZN(_06999_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15030_ (.A1(_06969_),
    .A2(_06998_),
    .B(_06999_),
    .ZN(_07000_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _15031_ (.A1(_06997_),
    .A2(_07000_),
    .ZN(_07001_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15032_ (.A1(_06971_),
    .A2(_06974_),
    .ZN(_07002_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _15033_ (.A1(_06958_),
    .A2(_06975_),
    .B(_07002_),
    .ZN(_07003_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _15034_ (.A1(_07001_),
    .A2(_07003_),
    .Z(_07004_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15035_ (.A1(_06983_),
    .A2(_07004_),
    .ZN(_07005_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15036_ (.A1(_06980_),
    .A2(_07005_),
    .B(_06979_),
    .ZN(_00562_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _15037_ (.A1(_06997_),
    .A2(_07000_),
    .Z(_07006_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15038_ (.A1(_07001_),
    .A2(_07003_),
    .B(_07006_),
    .ZN(_07007_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15039_ (.A1(_05969_),
    .A2(_06993_),
    .ZN(_07008_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15040_ (.A1(_05969_),
    .A2(_06993_),
    .ZN(_07009_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15041_ (.A1(_07008_),
    .A2(_06996_),
    .B(_07009_),
    .ZN(_07010_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _15042_ (.A1(_05014_),
    .A2(_05046_),
    .B(_04993_),
    .ZN(_07011_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _15043_ (.A1(_06994_),
    .A2(_06995_),
    .B(_07011_),
    .ZN(_07012_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _15044_ (.A1(_06986_),
    .A2(_06991_),
    .Z(_07013_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15045_ (.A1(_06984_),
    .A2(_06992_),
    .ZN(_07014_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _15046_ (.A1(_07013_),
    .A2(_07014_),
    .Z(_07015_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15047_ (.A1(_06989_),
    .A2(_06990_),
    .ZN(_07016_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15048_ (.A1(_06987_),
    .A2(_07016_),
    .ZN(_07017_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15049_ (.A1(_01769_),
    .A2(\channels.sample3[4] ),
    .ZN(_07018_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15050_ (.A1(_01760_),
    .A2(\channels.sample2[4] ),
    .ZN(_07019_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15051_ (.A1(_01746_),
    .A2(\channels.sample1[4] ),
    .ZN(_07020_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _15052_ (.A1(_07018_),
    .A2(_07019_),
    .A3(_07020_),
    .Z(_07021_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _15053_ (.A1(_07015_),
    .A2(_07017_),
    .A3(_07021_),
    .ZN(_07022_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _15054_ (.A1(\filters.low[5] ),
    .A2(_07022_),
    .Z(_07023_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _15055_ (.I(_07023_),
    .ZN(_07024_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _15056_ (.A1(_04992_),
    .A2(_07012_),
    .A3(_07024_),
    .Z(_07025_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _15057_ (.A1(_07010_),
    .A2(_07025_),
    .ZN(_07026_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _15058_ (.A1(_07010_),
    .A2(_07025_),
    .Z(_07027_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15059_ (.A1(_07026_),
    .A2(_07027_),
    .ZN(_07028_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15060_ (.I(_06981_),
    .Z(_07029_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _15061_ (.I(_07029_),
    .Z(_07030_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15062_ (.A1(_07007_),
    .A2(_07028_),
    .B(_07030_),
    .ZN(_07031_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15063_ (.A1(_07007_),
    .A2(_07028_),
    .B(_07031_),
    .ZN(_07032_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _15064_ (.I(_06982_),
    .Z(_07033_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15065_ (.A1(\filters.high[5] ),
    .A2(_07033_),
    .B(_06899_),
    .ZN(_07034_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15066_ (.A1(_07032_),
    .A2(_07034_),
    .ZN(_00563_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15067_ (.I(_07030_),
    .Z(_07035_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _15068_ (.A1(_07001_),
    .A2(_07003_),
    .B(_07027_),
    .C(_07006_),
    .ZN(_07036_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15069_ (.A1(_07026_),
    .A2(_07036_),
    .ZN(_07037_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _15070_ (.A1(_07017_),
    .A2(_07021_),
    .Z(_07038_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _15071_ (.A1(_07017_),
    .A2(_07021_),
    .Z(_07039_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15072_ (.A1(_07015_),
    .A2(_07038_),
    .B(_07039_),
    .ZN(_07040_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _15073_ (.A1(_07019_),
    .A2(_07020_),
    .Z(_07041_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _15074_ (.A1(_07019_),
    .A2(_07020_),
    .Z(_07042_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15075_ (.A1(_07018_),
    .A2(_07041_),
    .B(_07042_),
    .ZN(_07043_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15076_ (.A1(_01769_),
    .A2(\channels.sample3[5] ),
    .ZN(_07044_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15077_ (.A1(_01759_),
    .A2(\channels.sample2[5] ),
    .ZN(_07045_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15078_ (.A1(_01745_),
    .A2(\channels.sample1[5] ),
    .ZN(_07046_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _15079_ (.A1(_07045_),
    .A2(_07046_),
    .Z(_07047_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _15080_ (.A1(_07044_),
    .A2(_07047_),
    .Z(_07048_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _15081_ (.I(_07048_),
    .ZN(_07049_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _15082_ (.A1(_07043_),
    .A2(_07049_),
    .Z(_07050_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _15083_ (.A1(_07040_),
    .A2(_07050_),
    .Z(_07051_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _15084_ (.A1(\filters.low[6] ),
    .A2(_07051_),
    .Z(_07052_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _15085_ (.A1(net31),
    .A2(_05043_),
    .A3(_05048_),
    .ZN(_07053_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _15086_ (.A1(_07053_),
    .A2(_05421_),
    .Z(_07054_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _15087_ (.A1(_07052_),
    .A2(_07054_),
    .Z(_07055_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _15088_ (.A1(_04992_),
    .A2(_07012_),
    .ZN(_07056_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15089_ (.A1(_03310_),
    .A2(_07022_),
    .ZN(_07057_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _15090_ (.I(_07057_),
    .ZN(_07058_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _15091_ (.A1(_07056_),
    .A2(_07024_),
    .B(_07058_),
    .ZN(_07059_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _15092_ (.A1(_07055_),
    .A2(_07059_),
    .Z(_07060_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _15093_ (.A1(_07037_),
    .A2(_07060_),
    .Z(_07061_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _15094_ (.I(_06982_),
    .Z(_07062_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15095_ (.A1(\filters.high[6] ),
    .A2(_07062_),
    .B(_06775_),
    .ZN(_07063_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15096_ (.A1(_07035_),
    .A2(_07061_),
    .B(_07063_),
    .ZN(_00564_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15097_ (.I(_06913_),
    .Z(_07064_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _15098_ (.A1(_05417_),
    .A2(_05420_),
    .Z(_07065_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _15099_ (.A1(_07053_),
    .A2(_05421_),
    .B(_07065_),
    .ZN(_07066_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15100_ (.A1(_07043_),
    .A2(_07049_),
    .ZN(_07067_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15101_ (.A1(_07040_),
    .A2(_07050_),
    .ZN(_07068_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15102_ (.A1(_07067_),
    .A2(_07068_),
    .ZN(_07069_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15103_ (.A1(_01770_),
    .A2(_01927_),
    .A3(_07047_),
    .ZN(_07070_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15104_ (.A1(_07045_),
    .A2(_07046_),
    .B(_07070_),
    .ZN(_07071_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _15105_ (.I(_07071_),
    .ZN(_07072_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15106_ (.A1(_01769_),
    .A2(\channels.sample3[6] ),
    .ZN(_07073_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15107_ (.A1(_01760_),
    .A2(\channels.sample2[6] ),
    .ZN(_07074_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15108_ (.A1(_01746_),
    .A2(\channels.sample1[6] ),
    .ZN(_07075_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _15109_ (.A1(_07073_),
    .A2(_07074_),
    .A3(_07075_),
    .Z(_07076_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _15110_ (.A1(_07069_),
    .A2(_07072_),
    .A3(_07076_),
    .Z(_07077_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _15111_ (.A1(\filters.low[7] ),
    .A2(_07077_),
    .Z(_07078_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _15112_ (.A1(_05416_),
    .A2(_07066_),
    .A3(_07078_),
    .Z(_07079_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15113_ (.A1(_03329_),
    .A2(_07051_),
    .ZN(_07080_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _15114_ (.A1(_07052_),
    .A2(_07054_),
    .B(_07080_),
    .ZN(_07081_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _15115_ (.A1(_07079_),
    .A2(_07081_),
    .Z(_07082_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15116_ (.A1(_07055_),
    .A2(_07059_),
    .ZN(_07083_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15117_ (.A1(_07026_),
    .A2(_07036_),
    .A3(_07060_),
    .ZN(_07084_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _15118_ (.A1(_07083_),
    .A2(_07084_),
    .Z(_07085_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _15119_ (.I(_07029_),
    .Z(_07086_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15120_ (.A1(_07082_),
    .A2(_07085_),
    .B(_07086_),
    .ZN(_07087_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15121_ (.A1(_07082_),
    .A2(_07085_),
    .B(_07087_),
    .ZN(_07088_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15122_ (.I(_06186_),
    .Z(_07089_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _15123_ (.A1(_03343_),
    .A2(_07064_),
    .B(_07088_),
    .C(_07089_),
    .ZN(_00565_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _15124_ (.A1(_07055_),
    .A2(_07059_),
    .Z(_07090_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15125_ (.A1(_07079_),
    .A2(_07081_),
    .ZN(_07091_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15126_ (.A1(_07079_),
    .A2(_07081_),
    .ZN(_07092_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _15127_ (.A1(_07090_),
    .A2(_07091_),
    .B(_07092_),
    .ZN(_07093_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _15128_ (.A1(_07026_),
    .A2(_07036_),
    .A3(_07060_),
    .A4(_07082_),
    .ZN(_07094_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15129_ (.A1(_07093_),
    .A2(_07094_),
    .ZN(_07095_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15130_ (.A1(_05427_),
    .A2(_05428_),
    .ZN(_07096_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_4 _15131_ (.A1(_07053_),
    .A2(_05416_),
    .A3(_05421_),
    .B(_07096_),
    .ZN(_07097_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _15132_ (.A1(_05404_),
    .A2(_07097_),
    .ZN(_07098_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15133_ (.A1(_07072_),
    .A2(_07076_),
    .ZN(_07099_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15134_ (.A1(_07072_),
    .A2(_07076_),
    .ZN(_07100_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15135_ (.A1(_07069_),
    .A2(_07099_),
    .B(_07100_),
    .ZN(_07101_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _15136_ (.I(_07073_),
    .ZN(_07102_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15137_ (.A1(_07074_),
    .A2(_07075_),
    .ZN(_07103_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15138_ (.A1(_07074_),
    .A2(_07075_),
    .ZN(_07104_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _15139_ (.A1(_07102_),
    .A2(_07103_),
    .B(_07104_),
    .ZN(_07105_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15140_ (.A1(_01770_),
    .A2(\channels.sample3[7] ),
    .ZN(_07106_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15141_ (.A1(_01760_),
    .A2(\channels.sample2[7] ),
    .ZN(_07107_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15142_ (.A1(_01746_),
    .A2(\channels.sample1[7] ),
    .ZN(_07108_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _15143_ (.A1(_07107_),
    .A2(_07108_),
    .Z(_07109_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _15144_ (.A1(_07106_),
    .A2(_07109_),
    .Z(_07110_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _15145_ (.A1(_07101_),
    .A2(_07105_),
    .A3(_07110_),
    .ZN(_07111_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _15146_ (.A1(\filters.low[8] ),
    .A2(_07111_),
    .ZN(_07112_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _15147_ (.A1(_07098_),
    .A2(_07112_),
    .Z(_07113_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _15148_ (.A1(_05416_),
    .A2(_07066_),
    .ZN(_07114_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _15149_ (.A1(_03345_),
    .A2(_07077_),
    .Z(_07115_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _15150_ (.I(_07115_),
    .ZN(_07116_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _15151_ (.A1(_07114_),
    .A2(_07078_),
    .B(_07116_),
    .ZN(_07117_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _15152_ (.A1(_07113_),
    .A2(_07117_),
    .Z(_07118_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _15153_ (.A1(_07095_),
    .A2(_07118_),
    .Z(_07119_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15154_ (.A1(_06913_),
    .A2(_07119_),
    .ZN(_07120_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _15155_ (.A1(_03359_),
    .A2(_07064_),
    .B(_07120_),
    .C(_07089_),
    .ZN(_00566_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15156_ (.A1(_05379_),
    .A2(_05403_),
    .ZN(_07121_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _15157_ (.A1(_07121_),
    .A2(_07097_),
    .B(_05425_),
    .ZN(_07122_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _15158_ (.A1(_07105_),
    .A2(_07110_),
    .Z(_07123_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _15159_ (.A1(_07105_),
    .A2(_07110_),
    .Z(_07124_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15160_ (.A1(_07101_),
    .A2(_07123_),
    .B(_07124_),
    .ZN(_07125_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15161_ (.A1(_01771_),
    .A2(_01977_),
    .A3(_07109_),
    .ZN(_07126_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15162_ (.A1(_07107_),
    .A2(_07108_),
    .B(_07126_),
    .ZN(_07127_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _15163_ (.I(_07127_),
    .ZN(_07128_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15164_ (.A1(_01770_),
    .A2(\channels.sample3[8] ),
    .ZN(_07129_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15165_ (.A1(_01761_),
    .A2(\channels.sample2[8] ),
    .ZN(_07130_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15166_ (.A1(_01747_),
    .A2(\channels.sample1[8] ),
    .ZN(_07131_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _15167_ (.A1(_07129_),
    .A2(_07130_),
    .A3(_07131_),
    .Z(_07132_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _15168_ (.A1(_07125_),
    .A2(_07128_),
    .A3(_07132_),
    .Z(_07133_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _15169_ (.A1(\filters.low[9] ),
    .A2(_07133_),
    .ZN(_07134_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _15170_ (.A1(net56),
    .A2(_07122_),
    .A3(_07134_),
    .Z(_07135_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _15171_ (.I(_07112_),
    .ZN(_07136_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15172_ (.A1(_03360_),
    .A2(_07111_),
    .ZN(_07137_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _15173_ (.A1(_07098_),
    .A2(_07136_),
    .B(_07137_),
    .ZN(_07138_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _15174_ (.A1(_07135_),
    .A2(_07138_),
    .Z(_07139_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15175_ (.A1(_07113_),
    .A2(_07117_),
    .ZN(_07140_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15176_ (.A1(_07095_),
    .A2(_07118_),
    .B(_07140_),
    .ZN(_07141_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15177_ (.A1(_07139_),
    .A2(_07141_),
    .B(_07086_),
    .ZN(_07142_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15178_ (.A1(_07139_),
    .A2(_07141_),
    .B(_07142_),
    .ZN(_07143_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _15179_ (.A1(_03373_),
    .A2(_07064_),
    .B(_07143_),
    .C(_07089_),
    .ZN(_00567_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _15180_ (.A1(_07113_),
    .A2(_07117_),
    .ZN(_07144_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _15181_ (.A1(_07135_),
    .A2(_07138_),
    .ZN(_07145_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _15182_ (.A1(_07093_),
    .A2(_07094_),
    .B(_07144_),
    .C(_07145_),
    .ZN(_07146_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15183_ (.A1(_07135_),
    .A2(_07138_),
    .ZN(_07147_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _15184_ (.A1(_07113_),
    .A2(_07117_),
    .B1(_07135_),
    .B2(_07138_),
    .ZN(_07148_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _15185_ (.A1(_07147_),
    .A2(_07148_),
    .Z(_07149_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15186_ (.A1(_07128_),
    .A2(_07132_),
    .ZN(_07150_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15187_ (.A1(_07128_),
    .A2(_07132_),
    .ZN(_07151_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15188_ (.A1(_07125_),
    .A2(_07150_),
    .B(_07151_),
    .ZN(_07152_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _15189_ (.I(_07129_),
    .ZN(_07153_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15190_ (.A1(_07130_),
    .A2(_07131_),
    .ZN(_07154_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15191_ (.A1(_07130_),
    .A2(_07131_),
    .ZN(_07155_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15192_ (.A1(_07153_),
    .A2(_07154_),
    .B(_07155_),
    .ZN(_07156_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15193_ (.A1(_01771_),
    .A2(\channels.sample3[9] ),
    .ZN(_07157_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15194_ (.A1(_01761_),
    .A2(\channels.sample2[9] ),
    .ZN(_07158_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15195_ (.A1(_01747_),
    .A2(\channels.sample1[9] ),
    .ZN(_07159_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _15196_ (.A1(_07158_),
    .A2(_07159_),
    .Z(_07160_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _15197_ (.A1(_07157_),
    .A2(_07160_),
    .Z(_07161_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _15198_ (.A1(_07152_),
    .A2(_07156_),
    .A3(_07161_),
    .ZN(_07162_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _15199_ (.A1(\filters.low[10] ),
    .A2(_05532_),
    .A3(_07162_),
    .Z(_07163_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _15200_ (.I(_07163_),
    .ZN(_07164_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _15201_ (.A1(net56),
    .A2(_07122_),
    .Z(_07165_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _15202_ (.I(_07134_),
    .ZN(_07166_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15203_ (.A1(_03374_),
    .A2(_07133_),
    .ZN(_07167_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _15204_ (.A1(_07165_),
    .A2(_07166_),
    .B(_07167_),
    .ZN(_07168_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _15205_ (.A1(_07164_),
    .A2(_07168_),
    .Z(_07169_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15206_ (.A1(_07146_),
    .A2(_07149_),
    .B(_07169_),
    .ZN(_07170_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _15207_ (.A1(_07169_),
    .A2(_07146_),
    .A3(_07149_),
    .ZN(_07171_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15208_ (.A1(_06909_),
    .A2(_07171_),
    .ZN(_07172_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _15209_ (.A1(\filters.high[10] ),
    .A2(_06934_),
    .B1(_07170_),
    .B2(_07172_),
    .ZN(_07173_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15210_ (.A1(_06918_),
    .A2(_07173_),
    .ZN(_00568_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15211_ (.A1(_03394_),
    .A2(_07162_),
    .ZN(_07174_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15212_ (.A1(_03394_),
    .A2(_07162_),
    .ZN(_07175_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _15213_ (.A1(_05533_),
    .A2(_07174_),
    .B(_07175_),
    .ZN(_07176_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _15214_ (.A1(_07156_),
    .A2(_07161_),
    .Z(_07177_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _15215_ (.A1(_07156_),
    .A2(_07161_),
    .Z(_07178_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15216_ (.A1(_07152_),
    .A2(_07177_),
    .B(_07178_),
    .ZN(_07179_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15217_ (.A1(_01772_),
    .A2(_02029_),
    .A3(_07160_),
    .ZN(_07180_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15218_ (.A1(_07158_),
    .A2(_07159_),
    .B(_07180_),
    .ZN(_07181_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _15219_ (.I(_07181_),
    .ZN(_07182_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15220_ (.A1(_01771_),
    .A2(\channels.sample3[10] ),
    .ZN(_07183_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15221_ (.A1(_01762_),
    .A2(\channels.sample2[10] ),
    .ZN(_07184_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15222_ (.A1(_01748_),
    .A2(\channels.sample1[10] ),
    .ZN(_07185_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _15223_ (.A1(_07183_),
    .A2(_07184_),
    .A3(_07185_),
    .Z(_07186_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _15224_ (.A1(_07179_),
    .A2(_07182_),
    .A3(_07186_),
    .Z(_07187_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _15225_ (.A1(\filters.low[11] ),
    .A2(_07187_),
    .Z(_07188_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15226_ (.A1(_03411_),
    .A2(_07187_),
    .ZN(_07189_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15227_ (.A1(_07188_),
    .A2(_07189_),
    .ZN(_07190_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _15228_ (.A1(_07190_),
    .A2(_05646_),
    .ZN(_07191_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _15229_ (.A1(_07176_),
    .A2(_07191_),
    .ZN(_07192_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15230_ (.A1(_07164_),
    .A2(_07168_),
    .B(_07170_),
    .ZN(_07193_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15231_ (.A1(_07192_),
    .A2(_07193_),
    .B(_07086_),
    .ZN(_07194_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15232_ (.A1(_07192_),
    .A2(_07193_),
    .B(_07194_),
    .ZN(_07195_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _15233_ (.A1(_03410_),
    .A2(_07064_),
    .B(_07195_),
    .C(_07089_),
    .ZN(_00569_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _15234_ (.A1(_07176_),
    .A2(_07191_),
    .Z(_07196_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _15235_ (.A1(_07146_),
    .A2(_07149_),
    .B(_07196_),
    .C(_07169_),
    .ZN(_07197_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15236_ (.A1(_07164_),
    .A2(_07168_),
    .ZN(_07198_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15237_ (.A1(_07176_),
    .A2(_07191_),
    .ZN(_07199_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15238_ (.A1(_07176_),
    .A2(_07191_),
    .ZN(_07200_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _15239_ (.A1(_07198_),
    .A2(_07199_),
    .B(_07200_),
    .ZN(_07201_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15240_ (.A1(_07197_),
    .A2(_07201_),
    .ZN(_07202_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _15241_ (.I(_07202_),
    .ZN(_07203_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15242_ (.A1(_07182_),
    .A2(_07186_),
    .ZN(_07204_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15243_ (.A1(_07182_),
    .A2(_07186_),
    .ZN(_07205_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _15244_ (.A1(_07179_),
    .A2(_07204_),
    .B(_07205_),
    .ZN(_07206_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _15245_ (.I(_07183_),
    .ZN(_07207_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15246_ (.A1(_07184_),
    .A2(_07185_),
    .ZN(_07208_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15247_ (.A1(_07184_),
    .A2(_07185_),
    .ZN(_07209_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15248_ (.A1(_07207_),
    .A2(_07208_),
    .B(_07209_),
    .ZN(_07210_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15249_ (.A1(_01772_),
    .A2(\channels.sample3[11] ),
    .ZN(_07211_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15250_ (.A1(_01761_),
    .A2(\channels.sample2[11] ),
    .ZN(_07212_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15251_ (.A1(_01747_),
    .A2(\channels.sample1[11] ),
    .ZN(_07213_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _15252_ (.A1(_07212_),
    .A2(_07213_),
    .Z(_07214_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _15253_ (.A1(_07211_),
    .A2(_07214_),
    .Z(_07215_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _15254_ (.A1(_07206_),
    .A2(_07210_),
    .A3(_07215_),
    .ZN(_07216_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _15255_ (.A1(\filters.low[12] ),
    .A2(_07216_),
    .Z(_07217_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15256_ (.A1(_03422_),
    .A2(_07216_),
    .ZN(_07218_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _15257_ (.A1(_07217_),
    .A2(_07218_),
    .ZN(_07219_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15258_ (.A1(_05646_),
    .A2(_07190_),
    .B(_07188_),
    .ZN(_07220_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _15259_ (.A1(_05751_),
    .A2(_07219_),
    .A3(_07220_),
    .Z(_07221_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _15260_ (.A1(_07203_),
    .A2(_07221_),
    .Z(_07222_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15261_ (.I(_03721_),
    .Z(_07223_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15262_ (.A1(\filters.high[12] ),
    .A2(_07062_),
    .B(_07223_),
    .ZN(_07224_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15263_ (.A1(_07035_),
    .A2(_07222_),
    .B(_07224_),
    .ZN(_00570_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15264_ (.A1(_05751_),
    .A2(_07219_),
    .B(_07217_),
    .ZN(_07225_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15265_ (.A1(_01772_),
    .A2(_02056_),
    .A3(_07214_),
    .ZN(_07226_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _15266_ (.A1(_07212_),
    .A2(_07213_),
    .B(_07226_),
    .ZN(_07227_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _15267_ (.A1(_07210_),
    .A2(_07215_),
    .Z(_07228_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _15268_ (.A1(_07210_),
    .A2(_07215_),
    .Z(_07229_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _15269_ (.A1(_07206_),
    .A2(_07228_),
    .B(_07229_),
    .ZN(_07230_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _15270_ (.A1(_07227_),
    .A2(_07230_),
    .Z(_07231_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _15271_ (.A1(\filters.low[13] ),
    .A2(_07231_),
    .Z(_07232_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _15272_ (.I(_07232_),
    .ZN(_07233_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _15273_ (.A1(_05849_),
    .A2(_05851_),
    .A3(_07233_),
    .Z(_07234_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _15274_ (.A1(_07225_),
    .A2(_07234_),
    .ZN(_07235_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15275_ (.A1(_05752_),
    .A2(_07219_),
    .ZN(_07236_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _15276_ (.A1(_05751_),
    .A2(_07219_),
    .Z(_07237_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _15277_ (.A1(_07236_),
    .A2(_07237_),
    .A3(_07220_),
    .Z(_07238_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15278_ (.A1(_07202_),
    .A2(_07221_),
    .B(_07238_),
    .ZN(_07239_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _15279_ (.I(_07029_),
    .Z(_07240_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15280_ (.A1(_07235_),
    .A2(_07239_),
    .B(_07240_),
    .ZN(_07241_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15281_ (.A1(_07235_),
    .A2(_07239_),
    .B(_07241_),
    .ZN(_07242_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15282_ (.A1(\filters.high[13] ),
    .A2(_07033_),
    .B(_06899_),
    .ZN(_07243_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15283_ (.A1(_07242_),
    .A2(_07243_),
    .ZN(_00571_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _15284_ (.A1(_07227_),
    .A2(_07230_),
    .Z(_07244_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _15285_ (.A1(\filters.low[14] ),
    .A2(_07244_),
    .Z(_07245_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _15286_ (.A1(_05968_),
    .A2(_07245_),
    .Z(_07246_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15287_ (.A1(_03439_),
    .A2(_07231_),
    .ZN(_07247_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _15288_ (.I(_07247_),
    .ZN(_07248_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _15289_ (.A1(_05852_),
    .A2(_07233_),
    .B(_07248_),
    .ZN(_07249_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _15290_ (.A1(_07246_),
    .A2(_07249_),
    .Z(_07250_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15291_ (.A1(_07235_),
    .A2(_07221_),
    .ZN(_07251_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15292_ (.A1(_07217_),
    .A2(_07237_),
    .B(_07234_),
    .ZN(_07252_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15293_ (.A1(_07217_),
    .A2(_07237_),
    .A3(_07234_),
    .ZN(_07253_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _15294_ (.A1(_07238_),
    .A2(_07252_),
    .B(_07253_),
    .ZN(_07254_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15295_ (.A1(_07203_),
    .A2(_07251_),
    .B(_07254_),
    .ZN(_07255_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _15296_ (.A1(_07250_),
    .A2(_07255_),
    .Z(_07256_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15297_ (.A1(_07250_),
    .A2(_07255_),
    .B(_06982_),
    .ZN(_07257_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15298_ (.A1(_07256_),
    .A2(_07257_),
    .ZN(_07258_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15299_ (.A1(\filters.high[14] ),
    .A2(_06955_),
    .B(_07258_),
    .ZN(_07259_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15300_ (.A1(_06918_),
    .A2(_07259_),
    .ZN(_00572_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _15301_ (.A1(\filters.low[15] ),
    .A2(_06065_),
    .ZN(_07260_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15302_ (.A1(_05968_),
    .A2(_07245_),
    .ZN(_07261_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _15303_ (.A1(_03455_),
    .A2(_07244_),
    .B(_07261_),
    .ZN(_07262_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _15304_ (.A1(_07260_),
    .A2(_07262_),
    .Z(_07263_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _15305_ (.A1(_07260_),
    .A2(_07262_),
    .ZN(_07264_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15306_ (.A1(_07263_),
    .A2(_07264_),
    .ZN(_07265_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15307_ (.A1(_07246_),
    .A2(_07249_),
    .B(_07256_),
    .ZN(_07266_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15308_ (.A1(_07265_),
    .A2(_07266_),
    .B(_07086_),
    .ZN(_07267_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15309_ (.A1(_07265_),
    .A2(_07266_),
    .B(_07267_),
    .ZN(_07268_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _15310_ (.I(_06186_),
    .Z(_07269_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _15311_ (.A1(_03467_),
    .A2(_06910_),
    .B(_07268_),
    .C(_07269_),
    .ZN(_00573_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _15312_ (.A1(_07197_),
    .A2(_07201_),
    .B(_07251_),
    .ZN(_07270_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _15313_ (.A1(_07246_),
    .A2(_07249_),
    .ZN(_07271_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _15314_ (.A1(_07271_),
    .A2(_07263_),
    .A3(_07264_),
    .ZN(_07272_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _15315_ (.A1(_07271_),
    .A2(_07254_),
    .A3(_07263_),
    .A4(_07264_),
    .ZN(_07273_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15316_ (.A1(_07246_),
    .A2(_07249_),
    .ZN(_07274_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15317_ (.A1(_07260_),
    .A2(_07262_),
    .ZN(_07275_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _15318_ (.A1(_07274_),
    .A2(_07264_),
    .B(_07275_),
    .ZN(_07276_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _15319_ (.A1(_07270_),
    .A2(_07272_),
    .B(_07273_),
    .C(_07276_),
    .ZN(_07277_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15320_ (.A1(_03468_),
    .A2(_06065_),
    .ZN(_07278_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _15321_ (.A1(\filters.low[16] ),
    .A2(_06176_),
    .ZN(_07279_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _15322_ (.A1(_07278_),
    .A2(_07279_),
    .ZN(_07280_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _15323_ (.A1(_07277_),
    .A2(_07280_),
    .ZN(_07281_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15324_ (.A1(\filters.high[16] ),
    .A2(_07062_),
    .B(_07223_),
    .ZN(_07282_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15325_ (.A1(_07035_),
    .A2(_07281_),
    .B(_07282_),
    .ZN(_00574_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _15326_ (.A1(\filters.low[16] ),
    .A2(_06287_),
    .Z(_07283_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _15327_ (.A1(\filters.low[17] ),
    .A2(_06293_),
    .A3(_07283_),
    .ZN(_07284_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15328_ (.A1(_07278_),
    .A2(_07279_),
    .ZN(_07285_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15329_ (.A1(_07277_),
    .A2(_07280_),
    .B(_07285_),
    .ZN(_07286_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _15330_ (.A1(_07284_),
    .A2(_07286_),
    .ZN(_07287_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15331_ (.A1(_06919_),
    .A2(_07287_),
    .ZN(_07288_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15332_ (.A1(\filters.high[17] ),
    .A2(_07033_),
    .B(_06899_),
    .ZN(_07289_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15333_ (.A1(_07288_),
    .A2(_07289_),
    .ZN(_00575_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15334_ (.A1(\filters.high[18] ),
    .A2(_06955_),
    .ZN(_07290_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15335_ (.A1(\filters.low[17] ),
    .A2(_06293_),
    .ZN(_07291_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _15336_ (.A1(\filters.low[18] ),
    .A2(_06396_),
    .Z(_07292_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _15337_ (.A1(_07291_),
    .A2(_07292_),
    .Z(_07293_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _15338_ (.A1(_07280_),
    .A2(_07284_),
    .Z(_07294_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _15339_ (.I(\filters.low[17] ),
    .Z(_07295_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _15340_ (.A1(_07295_),
    .A2(_06294_),
    .Z(_07296_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15341_ (.A1(_07283_),
    .A2(_07296_),
    .ZN(_07297_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15342_ (.A1(_07283_),
    .A2(_07296_),
    .B(_07285_),
    .ZN(_07298_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _15343_ (.A1(_07297_),
    .A2(_07298_),
    .ZN(_07299_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15344_ (.A1(_07277_),
    .A2(_07294_),
    .B(_07299_),
    .ZN(_07300_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _15345_ (.A1(_07293_),
    .A2(_07300_),
    .ZN(_07301_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15346_ (.A1(_06983_),
    .A2(_07301_),
    .ZN(_07302_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15347_ (.A1(_07290_),
    .A2(_07302_),
    .B(_06979_),
    .ZN(_00576_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _15348_ (.A1(\filters.low[18] ),
    .A2(_06396_),
    .Z(_07303_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _15349_ (.A1(\filters.low[19] ),
    .A2(_06498_),
    .Z(_07304_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _15350_ (.A1(_07303_),
    .A2(_07304_),
    .ZN(_07305_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15351_ (.A1(_07295_),
    .A2(_06294_),
    .A3(_07292_),
    .ZN(_07306_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _15352_ (.A1(_07295_),
    .A2(_06294_),
    .B(_07292_),
    .ZN(_07307_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15353_ (.A1(_07306_),
    .A2(_07300_),
    .B(_07307_),
    .ZN(_07308_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _15354_ (.A1(_07305_),
    .A2(_07308_),
    .ZN(_07309_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15355_ (.I(_07029_),
    .Z(_07310_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15356_ (.A1(\filters.high[19] ),
    .A2(_07310_),
    .B(_07223_),
    .ZN(_07311_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15357_ (.A1(_07035_),
    .A2(_07309_),
    .B(_07311_),
    .ZN(_00577_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15358_ (.I(_07030_),
    .Z(_07312_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15359_ (.A1(\filters.low[19] ),
    .A2(_06499_),
    .ZN(_07313_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _15360_ (.A1(\filters.low[20] ),
    .A2(_06599_),
    .ZN(_07314_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _15361_ (.A1(_07313_),
    .A2(_07314_),
    .Z(_07315_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _15362_ (.A1(_07293_),
    .A2(_07305_),
    .Z(_07316_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _15363_ (.A1(_07293_),
    .A2(_07294_),
    .A3(_07305_),
    .Z(_07317_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15364_ (.A1(_07303_),
    .A2(_07304_),
    .ZN(_07318_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15365_ (.A1(_07303_),
    .A2(_07304_),
    .ZN(_07319_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _15366_ (.A1(_07307_),
    .A2(_07318_),
    .B(_07319_),
    .ZN(_07320_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _15367_ (.A1(_07299_),
    .A2(_07316_),
    .B1(_07317_),
    .B2(_07277_),
    .C(_07320_),
    .ZN(_07321_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _15368_ (.A1(_07315_),
    .A2(_07321_),
    .ZN(_07322_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15369_ (.A1(\filters.high[20] ),
    .A2(_07310_),
    .B(_07223_),
    .ZN(_07323_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15370_ (.A1(_07312_),
    .A2(_07322_),
    .B(_07323_),
    .ZN(_00578_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15371_ (.A1(_07313_),
    .A2(_07314_),
    .ZN(_07324_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15372_ (.A1(_07315_),
    .A2(_07321_),
    .ZN(_07325_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _15373_ (.A1(_07324_),
    .A2(_07325_),
    .Z(_07326_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15374_ (.I(\filters.low[21] ),
    .Z(_07327_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15375_ (.A1(\filters.low[20] ),
    .A2(_06599_),
    .ZN(_07328_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _15376_ (.A1(_07327_),
    .A2(_06754_),
    .A3(_07328_),
    .ZN(_07329_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15377_ (.A1(_07326_),
    .A2(_07329_),
    .B(_07240_),
    .ZN(_07330_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15378_ (.A1(_07326_),
    .A2(_07329_),
    .B(_07330_),
    .ZN(_07331_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15379_ (.I(_03733_),
    .Z(_07332_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _15380_ (.I(_07332_),
    .Z(_07333_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15381_ (.A1(\filters.high[21] ),
    .A2(_07033_),
    .B(_07333_),
    .ZN(_07334_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15382_ (.A1(_07331_),
    .A2(_07334_),
    .ZN(_00579_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15383_ (.A1(\filters.high[22] ),
    .A2(_06919_),
    .ZN(_07335_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _15384_ (.A1(_07315_),
    .A2(_07329_),
    .Z(_07336_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _15385_ (.A1(_07327_),
    .A2(_06836_),
    .ZN(_07337_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15386_ (.A1(_07328_),
    .A2(_07337_),
    .ZN(_07338_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15387_ (.A1(_07328_),
    .A2(_07337_),
    .ZN(_07339_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _15388_ (.A1(_07324_),
    .A2(_07338_),
    .B(_07339_),
    .ZN(_07340_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15389_ (.A1(_07321_),
    .A2(_07336_),
    .B(_07340_),
    .ZN(_07341_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _15390_ (.I(_07341_),
    .ZN(_07342_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15391_ (.A1(_07327_),
    .A2(_06716_),
    .ZN(_07343_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _15392_ (.A1(\filters.low[22] ),
    .A2(_06754_),
    .Z(_07344_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _15393_ (.A1(_07343_),
    .A2(_07344_),
    .ZN(_07345_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _15394_ (.A1(_07342_),
    .A2(_07345_),
    .Z(_07346_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15395_ (.A1(_07062_),
    .A2(_07346_),
    .ZN(_07347_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15396_ (.A1(_07335_),
    .A2(_07347_),
    .B(_06979_),
    .ZN(_00580_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _15397_ (.I(_07343_),
    .ZN(_07348_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15398_ (.A1(_07348_),
    .A2(_07344_),
    .ZN(_07349_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15399_ (.A1(_07342_),
    .A2(_07345_),
    .B(_07349_),
    .ZN(_07350_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15400_ (.A1(\filters.low[22] ),
    .A2(_06836_),
    .ZN(_07351_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _15401_ (.A1(\filters.low[23] ),
    .A2(_06701_),
    .Z(_07352_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _15402_ (.A1(_07351_),
    .A2(_07352_),
    .ZN(_07353_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _15403_ (.A1(_07350_),
    .A2(_07353_),
    .Z(_07354_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _15404_ (.I(_02100_),
    .Z(_07355_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _15405_ (.I(_07355_),
    .Z(_07356_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15406_ (.A1(\filters.high[23] ),
    .A2(_07310_),
    .B(_07356_),
    .ZN(_07357_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15407_ (.A1(_07312_),
    .A2(_07354_),
    .B(_07357_),
    .ZN(_00581_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _15408_ (.A1(_07345_),
    .A2(_07353_),
    .Z(_07358_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _15409_ (.A1(_07336_),
    .A2(_07345_),
    .A3(_07353_),
    .Z(_07359_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _15410_ (.I(_07351_),
    .ZN(_07360_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _15411_ (.A1(_06822_),
    .A2(_07348_),
    .A3(_07344_),
    .B1(_07352_),
    .B2(_07360_),
    .ZN(_07361_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _15412_ (.A1(_07340_),
    .A2(_07358_),
    .B1(_07359_),
    .B2(_07321_),
    .C(_07361_),
    .ZN(_07362_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _15413_ (.I(\filters.low[24] ),
    .Z(_07363_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _15414_ (.A1(_07363_),
    .A2(_06852_),
    .Z(_07364_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _15415_ (.A1(\filters.low[23] ),
    .A2(_06862_),
    .Z(_07365_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _15416_ (.I0(_07364_),
    .I1(_07363_),
    .S(_07365_),
    .Z(_07366_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _15417_ (.A1(_07362_),
    .A2(_07366_),
    .Z(_07367_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15418_ (.A1(\filters.high[24] ),
    .A2(_07310_),
    .B(_07356_),
    .ZN(_07368_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15419_ (.A1(_07312_),
    .A2(_07367_),
    .B(_07368_),
    .ZN(_00582_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _15420_ (.I(\filters.high[25] ),
    .ZN(_07369_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _15421_ (.A1(_07365_),
    .A2(_07364_),
    .ZN(_07370_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _15422_ (.A1(_06837_),
    .A2(_07365_),
    .B(_07362_),
    .C(_07370_),
    .ZN(_07371_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15423_ (.I(\filters.low[25] ),
    .Z(_07372_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _15424_ (.I(_07372_),
    .Z(_07373_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _15425_ (.A1(_07363_),
    .A2(_06862_),
    .ZN(_07374_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _15426_ (.A1(_07372_),
    .A2(_06852_),
    .Z(_07375_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _15427_ (.I(_07375_),
    .ZN(_07376_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15428_ (.A1(_07374_),
    .A2(_07376_),
    .ZN(_07377_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15429_ (.A1(_07373_),
    .A2(_07374_),
    .B(_07377_),
    .ZN(_07378_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15430_ (.A1(_07370_),
    .A2(_07371_),
    .B(_07378_),
    .ZN(_07379_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _15431_ (.A1(_07370_),
    .A2(_07371_),
    .A3(_07378_),
    .ZN(_07380_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15432_ (.A1(_06934_),
    .A2(_07380_),
    .ZN(_07381_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _15433_ (.A1(_07369_),
    .A2(_06910_),
    .B1(_07379_),
    .B2(_07381_),
    .C(_06917_),
    .ZN(_00583_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15434_ (.I(_01932_),
    .Z(_07382_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15435_ (.I(\filters.low[26] ),
    .Z(_07383_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _15436_ (.A1(\filters.low[26] ),
    .A2(_06852_),
    .Z(_07384_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15437_ (.A1(_07372_),
    .A2(_06765_),
    .ZN(_07385_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _15438_ (.I0(_07383_),
    .I1(_07384_),
    .S(_07385_),
    .Z(_07386_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _15439_ (.I0(_07372_),
    .I1(_07375_),
    .S(_07374_),
    .Z(_07387_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15440_ (.A1(_07366_),
    .A2(_07387_),
    .ZN(_07388_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _15441_ (.A1(_07373_),
    .A2(_07370_),
    .B1(_07376_),
    .B2(_07374_),
    .ZN(_07389_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15442_ (.A1(net36),
    .A2(_07388_),
    .B(_07389_),
    .ZN(_07390_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15443_ (.A1(_07386_),
    .A2(_07390_),
    .ZN(_07391_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15444_ (.A1(_07386_),
    .A2(_07390_),
    .ZN(_07392_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15445_ (.A1(_06909_),
    .A2(_07392_),
    .ZN(_07393_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _15446_ (.A1(\filters.high[26] ),
    .A2(_06934_),
    .B1(_07391_),
    .B2(_07393_),
    .ZN(_07394_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15447_ (.A1(_07382_),
    .A2(_07394_),
    .ZN(_00584_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _15448_ (.I(\filters.low[27] ),
    .Z(_07395_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _15449_ (.A1(\filters.low[27] ),
    .A2(_06862_),
    .Z(_07396_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15450_ (.A1(_07383_),
    .A2(_06734_),
    .ZN(_07397_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _15451_ (.I0(_07395_),
    .I1(_07396_),
    .S(_07397_),
    .Z(_07398_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _15452_ (.A1(_07373_),
    .A2(_06767_),
    .B(_07384_),
    .ZN(_07399_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15453_ (.A1(_07386_),
    .A2(_07390_),
    .B(_07399_),
    .ZN(_07400_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15454_ (.A1(_07398_),
    .A2(_07400_),
    .B(_07240_),
    .ZN(_07401_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15455_ (.A1(_07398_),
    .A2(_07400_),
    .B(_07401_),
    .ZN(_07402_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15456_ (.A1(\filters.high[27] ),
    .A2(_06983_),
    .B(_07333_),
    .ZN(_07403_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15457_ (.A1(_07402_),
    .A2(_07403_),
    .ZN(_00585_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15458_ (.A1(_07386_),
    .A2(_07398_),
    .ZN(_07404_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _15459_ (.A1(_07388_),
    .A2(_07404_),
    .Z(_07405_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15460_ (.A1(_07383_),
    .A2(_06767_),
    .B(_07396_),
    .ZN(_07406_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _15461_ (.A1(_07395_),
    .A2(_07399_),
    .B(_07406_),
    .ZN(_07407_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _15462_ (.A1(_07389_),
    .A2(_07404_),
    .B1(_07405_),
    .B2(_07362_),
    .C(_07407_),
    .ZN(_07408_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _15463_ (.A1(_07395_),
    .A2(_06766_),
    .Z(_07409_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _15464_ (.A1(\filters.low[28] ),
    .A2(_06717_),
    .Z(_07410_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _15465_ (.A1(_07409_),
    .A2(_07410_),
    .ZN(_07411_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _15466_ (.A1(_06875_),
    .A2(_07409_),
    .B(_07411_),
    .ZN(_07412_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _15467_ (.A1(_07408_),
    .A2(_07412_),
    .ZN(_07413_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15468_ (.A1(\filters.high[28] ),
    .A2(_07030_),
    .B(_07356_),
    .ZN(_07414_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15469_ (.A1(_07312_),
    .A2(_07413_),
    .B(_07414_),
    .ZN(_00586_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _15470_ (.A1(\filters.low[28] ),
    .A2(_06766_),
    .Z(_07415_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _15471_ (.I(\filters.low[29] ),
    .Z(_07416_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _15472_ (.A1(_07416_),
    .A2(_06717_),
    .Z(_07417_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _15473_ (.A1(_07415_),
    .A2(_07417_),
    .ZN(_07418_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _15474_ (.A1(_06882_),
    .A2(_07415_),
    .B(_07418_),
    .ZN(_07419_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15475_ (.A1(_07408_),
    .A2(_07412_),
    .B(_07411_),
    .ZN(_07420_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15476_ (.A1(_07419_),
    .A2(_07420_),
    .B(_07240_),
    .ZN(_07421_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15477_ (.A1(_07419_),
    .A2(_07420_),
    .B(_07421_),
    .ZN(_07422_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15478_ (.A1(\filters.high[29] ),
    .A2(_06983_),
    .B(_07333_),
    .ZN(_07423_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15479_ (.A1(_07422_),
    .A2(_07423_),
    .ZN(_00587_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15480_ (.A1(\filters.high[30] ),
    .A2(_06919_),
    .ZN(_07424_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _15481_ (.A1(_07412_),
    .A2(_07419_),
    .Z(_07425_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _15482_ (.A1(_07416_),
    .A2(_07411_),
    .B1(_07425_),
    .B2(_07408_),
    .C(_07418_),
    .ZN(_07426_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15483_ (.A1(_06891_),
    .A2(_06767_),
    .ZN(_07427_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _15484_ (.I(_07427_),
    .ZN(_07428_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15485_ (.A1(_06891_),
    .A2(_06719_),
    .ZN(_07429_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _15486_ (.A1(_07416_),
    .A2(_06768_),
    .B(_07429_),
    .C(_07428_),
    .ZN(_07430_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15487_ (.A1(_07416_),
    .A2(_07428_),
    .B(_07430_),
    .ZN(_07431_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _15488_ (.I(_07431_),
    .ZN(_07432_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15489_ (.A1(net67),
    .A2(_07432_),
    .B(_06952_),
    .ZN(_07433_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15490_ (.A1(_07426_),
    .A2(_07432_),
    .B(_07433_),
    .ZN(_07434_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15491_ (.I(_06978_),
    .Z(_07435_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15492_ (.A1(_07424_),
    .A2(_07434_),
    .B(_07435_),
    .ZN(_00588_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _15493_ (.I(\filters.high[31] ),
    .ZN(_07436_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _15494_ (.A1(_07426_),
    .A2(_07432_),
    .ZN(_07437_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _15495_ (.A1(_07430_),
    .A2(_07437_),
    .Z(_07438_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _15496_ (.A1(\filters.low[31] ),
    .A2(_07428_),
    .Z(_07439_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _15497_ (.I(_07439_),
    .ZN(_07440_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _15498_ (.A1(_07438_),
    .A2(_07440_),
    .Z(_07441_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15499_ (.A1(_07438_),
    .A2(_07440_),
    .B(_06913_),
    .ZN(_07442_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _15500_ (.A1(_07436_),
    .A2(_06910_),
    .B1(_07441_),
    .B2(_07442_),
    .C(_06917_),
    .ZN(_00589_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _15501_ (.I(_03202_),
    .Z(_07443_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _15502_ (.A1(\filters.mode_vol[7] ),
    .A2(_01773_),
    .B(_03214_),
    .C(_03215_),
    .ZN(_07444_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_4 _15503_ (.A1(_01748_),
    .A2(_03428_),
    .B1(_03476_),
    .B2(_01762_),
    .C1(_07443_),
    .C2(_03237_),
    .ZN(_07445_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _15504_ (.A1(_07443_),
    .A2(_07444_),
    .B(_07445_),
    .C(_03729_),
    .ZN(_07446_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15505_ (.I(_07446_),
    .Z(_07447_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15506_ (.I(_07447_),
    .Z(_07448_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _15507_ (.A1(_03194_),
    .A2(_04189_),
    .B(_07446_),
    .ZN(_07449_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15508_ (.I(_07449_),
    .Z(_07450_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15509_ (.I(_07450_),
    .Z(_07451_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _15510_ (.A1(_03202_),
    .A2(_03204_),
    .A3(_03215_),
    .ZN(_07452_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15511_ (.I(_07452_),
    .Z(_07453_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15512_ (.A1(\channels.sample3[0] ),
    .A2(_07453_),
    .ZN(_07454_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _15513_ (.A1(_03263_),
    .A2(_07453_),
    .B(_07454_),
    .C(_03219_),
    .ZN(_07455_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _15514_ (.A1(\channels.sample2[0] ),
    .A2(_06066_),
    .B(_07455_),
    .C(_03344_),
    .ZN(_07456_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15515_ (.A1(\channels.sample1[0] ),
    .A2(_03400_),
    .ZN(_07457_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _15516_ (.A1(_07456_),
    .A2(_07457_),
    .ZN(_07458_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _15517_ (.A1(\filters.sample_buff[0] ),
    .A2(_07458_),
    .Z(_07459_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _15518_ (.A1(\filters.sample_buff[0] ),
    .A2(_07448_),
    .B1(_07451_),
    .B2(_07459_),
    .ZN(_07460_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15519_ (.A1(_07382_),
    .A2(_07460_),
    .ZN(_00590_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15520_ (.I(_07446_),
    .Z(_07461_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _15521_ (.A1(\filters.sample_buff[0] ),
    .A2(_07458_),
    .Z(_07462_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _15522_ (.I(_07452_),
    .Z(_07463_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15523_ (.A1(\channels.sample3[1] ),
    .A2(_07452_),
    .ZN(_07464_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _15524_ (.A1(_03264_),
    .A2(_07463_),
    .B(_07464_),
    .C(_03218_),
    .ZN(_07465_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _15525_ (.A1(\channels.sample2[1] ),
    .A2(_03219_),
    .B(_07465_),
    .C(_03229_),
    .ZN(_07466_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15526_ (.A1(\channels.sample1[1] ),
    .A2(_03335_),
    .ZN(_07467_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _15527_ (.A1(_07466_),
    .A2(_07467_),
    .ZN(_07468_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _15528_ (.A1(\filters.sample_buff[1] ),
    .A2(_07468_),
    .Z(_07469_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _15529_ (.A1(_07462_),
    .A2(_07469_),
    .Z(_07470_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _15530_ (.A1(\filters.sample_buff[1] ),
    .A2(_07461_),
    .B1(_07451_),
    .B2(_07470_),
    .ZN(_07471_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15531_ (.A1(_07382_),
    .A2(_07471_),
    .ZN(_00591_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15532_ (.A1(\filters.sample_buff[1] ),
    .A2(_07468_),
    .ZN(_07472_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15533_ (.A1(_07462_),
    .A2(_07469_),
    .ZN(_07473_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15534_ (.A1(\channels.sample3[2] ),
    .A2(_07463_),
    .ZN(_07474_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _15535_ (.A1(_03281_),
    .A2(_07463_),
    .B(_07474_),
    .C(_03375_),
    .ZN(_07475_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _15536_ (.A1(\channels.sample2[2] ),
    .A2(_03346_),
    .B(_07475_),
    .C(_03229_),
    .ZN(_07476_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15537_ (.A1(\channels.sample1[2] ),
    .A2(_03335_),
    .ZN(_07477_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _15538_ (.A1(_07476_),
    .A2(_07477_),
    .ZN(_07478_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _15539_ (.A1(\filters.sample_buff[2] ),
    .A2(_07478_),
    .ZN(_07479_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _15540_ (.A1(_07472_),
    .A2(_07473_),
    .B(_07479_),
    .ZN(_07480_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _15541_ (.A1(_07472_),
    .A2(_07473_),
    .A3(_07479_),
    .Z(_07481_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15542_ (.A1(_07480_),
    .A2(_07481_),
    .ZN(_07482_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _15543_ (.A1(\filters.sample_buff[2] ),
    .A2(_07461_),
    .B1(_07451_),
    .B2(_07482_),
    .ZN(_07483_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15544_ (.A1(_07382_),
    .A2(_07483_),
    .ZN(_00592_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _15545_ (.I(_07446_),
    .Z(_07484_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15546_ (.A1(\filters.sample_buff[3] ),
    .A2(_07484_),
    .ZN(_07485_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15547_ (.I(_07449_),
    .Z(_07486_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _15548_ (.A1(\filters.sample_buff[2] ),
    .A2(_07478_),
    .Z(_07487_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _15549_ (.I(_07463_),
    .Z(_07488_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15550_ (.A1(\channels.sample3[3] ),
    .A2(_07453_),
    .ZN(_07489_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _15551_ (.A1(_03297_),
    .A2(_07488_),
    .B(_07489_),
    .C(_03376_),
    .ZN(_07490_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _15552_ (.A1(\channels.sample2[3] ),
    .A2(_03220_),
    .B(_07490_),
    .C(_03344_),
    .ZN(_07491_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15553_ (.A1(\channels.sample1[3] ),
    .A2(_03400_),
    .ZN(_07492_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _15554_ (.A1(_07491_),
    .A2(_07492_),
    .ZN(_07493_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _15555_ (.A1(\filters.sample_buff[3] ),
    .A2(_07493_),
    .Z(_07494_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _15556_ (.A1(_07487_),
    .A2(_07480_),
    .A3(_07494_),
    .Z(_07495_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _15557_ (.A1(_07487_),
    .A2(_07480_),
    .B(_07494_),
    .ZN(_07496_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15558_ (.A1(_07486_),
    .A2(_07495_),
    .A3(_07496_),
    .ZN(_07497_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15559_ (.A1(_07485_),
    .A2(_07497_),
    .B(_07435_),
    .ZN(_00593_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15560_ (.I(_01932_),
    .Z(_07498_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15561_ (.A1(\filters.sample_buff[3] ),
    .A2(_07493_),
    .ZN(_07499_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15562_ (.A1(\channels.sample3[4] ),
    .A2(_07453_),
    .ZN(_07500_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _15563_ (.A1(_03309_),
    .A2(_07488_),
    .B(_07500_),
    .C(_06066_),
    .ZN(_07501_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _15564_ (.A1(\channels.sample2[4] ),
    .A2(_03377_),
    .B(_07501_),
    .C(_03230_),
    .ZN(_07502_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15565_ (.A1(\channels.sample1[4] ),
    .A2(_03400_),
    .ZN(_07503_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _15566_ (.A1(_07502_),
    .A2(_07503_),
    .ZN(_07504_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _15567_ (.A1(\filters.sample_buff[4] ),
    .A2(_07504_),
    .Z(_07505_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _15568_ (.I(_07505_),
    .ZN(_07506_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _15569_ (.A1(_07499_),
    .A2(_07496_),
    .B(_07506_),
    .ZN(_07507_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _15570_ (.A1(_07499_),
    .A2(_07496_),
    .A3(_07506_),
    .Z(_07508_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15571_ (.A1(_07507_),
    .A2(_07508_),
    .ZN(_07509_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _15572_ (.A1(\filters.sample_buff[4] ),
    .A2(_07461_),
    .B1(_07451_),
    .B2(_07509_),
    .ZN(_07510_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15573_ (.A1(_07498_),
    .A2(_07510_),
    .ZN(_00594_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15574_ (.A1(\filters.sample_buff[5] ),
    .A2(_07484_),
    .ZN(_07511_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _15575_ (.A1(\filters.sample_buff[4] ),
    .A2(_07504_),
    .Z(_07512_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15576_ (.I(_07488_),
    .Z(_07513_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15577_ (.A1(_01927_),
    .A2(_07488_),
    .ZN(_07514_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _15578_ (.A1(_03326_),
    .A2(_07513_),
    .B(_07514_),
    .C(_06067_),
    .ZN(_07515_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _15579_ (.A1(\channels.sample2[5] ),
    .A2(_03378_),
    .B(_07515_),
    .C(_03231_),
    .ZN(_07516_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15580_ (.A1(\channels.sample1[5] ),
    .A2(_03401_),
    .ZN(_07517_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _15581_ (.A1(_07516_),
    .A2(_07517_),
    .ZN(_07518_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _15582_ (.A1(\filters.sample_buff[5] ),
    .A2(_07518_),
    .Z(_07519_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _15583_ (.A1(_07512_),
    .A2(_07507_),
    .A3(_07519_),
    .Z(_07520_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _15584_ (.A1(_07512_),
    .A2(_07507_),
    .B(_07519_),
    .ZN(_07521_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15585_ (.A1(_07486_),
    .A2(_07520_),
    .A3(_07521_),
    .ZN(_07522_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15586_ (.A1(_07511_),
    .A2(_07522_),
    .B(_07435_),
    .ZN(_00595_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15587_ (.I(_07449_),
    .Z(_07523_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15588_ (.A1(\filters.sample_buff[5] ),
    .A2(_07518_),
    .ZN(_07524_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15589_ (.A1(\channels.sample3[6] ),
    .A2(_07513_),
    .ZN(_07525_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _15590_ (.A1(_03342_),
    .A2(_07513_),
    .B(_07525_),
    .C(_06177_),
    .ZN(_07526_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _15591_ (.A1(\channels.sample2[6] ),
    .A2(_06397_),
    .B(_07526_),
    .C(_03231_),
    .ZN(_07527_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15592_ (.A1(\channels.sample1[6] ),
    .A2(_03401_),
    .ZN(_07528_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _15593_ (.A1(_07527_),
    .A2(_07528_),
    .ZN(_07529_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _15594_ (.A1(\filters.sample_buff[6] ),
    .A2(_07529_),
    .Z(_07530_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _15595_ (.I(_07530_),
    .ZN(_07531_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _15596_ (.A1(_07524_),
    .A2(_07521_),
    .B(_07531_),
    .ZN(_07532_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _15597_ (.A1(_07524_),
    .A2(_07521_),
    .A3(_07531_),
    .Z(_07533_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15598_ (.A1(_07532_),
    .A2(_07533_),
    .ZN(_07534_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _15599_ (.A1(\filters.sample_buff[6] ),
    .A2(_07461_),
    .B1(_07523_),
    .B2(_07534_),
    .ZN(_07535_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15600_ (.A1(_07498_),
    .A2(_07535_),
    .ZN(_00596_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15601_ (.A1(\filters.sample_buff[7] ),
    .A2(_07484_),
    .ZN(_07536_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _15602_ (.A1(\filters.sample_buff[6] ),
    .A2(_07529_),
    .Z(_07537_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15603_ (.I(_07513_),
    .Z(_07538_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15604_ (.A1(_01977_),
    .A2(_07538_),
    .ZN(_07539_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _15605_ (.A1(_03358_),
    .A2(_07538_),
    .B(_07539_),
    .C(_06710_),
    .ZN(_07540_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _15606_ (.A1(\channels.sample2[7] ),
    .A2(_03395_),
    .B(_07540_),
    .C(_03232_),
    .ZN(_07541_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15607_ (.A1(\channels.sample1[7] ),
    .A2(_03427_),
    .ZN(_07542_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _15608_ (.A1(_07541_),
    .A2(_07542_),
    .ZN(_07543_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _15609_ (.A1(\filters.sample_buff[7] ),
    .A2(_07543_),
    .Z(_07544_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _15610_ (.A1(_07537_),
    .A2(_07532_),
    .A3(_07544_),
    .Z(_07545_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _15611_ (.A1(_07537_),
    .A2(_07532_),
    .B(_07544_),
    .ZN(_07546_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15612_ (.A1(_07486_),
    .A2(_07545_),
    .A3(_07546_),
    .ZN(_07547_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15613_ (.A1(_07536_),
    .A2(_07547_),
    .B(_07435_),
    .ZN(_00597_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15614_ (.A1(\filters.sample_buff[7] ),
    .A2(_07543_),
    .ZN(_07548_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15615_ (.I(_07538_),
    .Z(_07549_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15616_ (.A1(\channels.sample3[8] ),
    .A2(_07538_),
    .ZN(_07550_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _15617_ (.A1(_03372_),
    .A2(_07549_),
    .B(_07550_),
    .C(_03395_),
    .ZN(_07551_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _15618_ (.A1(\channels.sample2[8] ),
    .A2(_03223_),
    .B(_07551_),
    .C(_03232_),
    .ZN(_07552_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15619_ (.A1(\channels.sample1[8] ),
    .A2(_03427_),
    .ZN(_07553_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _15620_ (.A1(_07552_),
    .A2(_07553_),
    .ZN(_07554_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _15621_ (.A1(\filters.sample_buff[8] ),
    .A2(_07554_),
    .Z(_07555_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _15622_ (.I(_07555_),
    .ZN(_07556_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _15623_ (.A1(_07548_),
    .A2(_07546_),
    .B(_07556_),
    .ZN(_07557_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _15624_ (.A1(_07548_),
    .A2(_07546_),
    .A3(_07556_),
    .Z(_07558_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15625_ (.A1(_07557_),
    .A2(_07558_),
    .ZN(_07559_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _15626_ (.A1(\filters.sample_buff[8] ),
    .A2(_07447_),
    .B1(_07523_),
    .B2(_07559_),
    .ZN(_07560_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15627_ (.A1(_07498_),
    .A2(_07560_),
    .ZN(_00598_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15628_ (.A1(\filters.sample_buff[9] ),
    .A2(_07448_),
    .ZN(_07561_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _15629_ (.A1(\filters.sample_buff[8] ),
    .A2(_07554_),
    .Z(_07562_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15630_ (.I(_07549_),
    .Z(_07563_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15631_ (.A1(_02029_),
    .A2(_07549_),
    .ZN(_07564_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _15632_ (.A1(_03391_),
    .A2(_07563_),
    .B(_07564_),
    .C(_03223_),
    .ZN(_07565_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _15633_ (.A1(\channels.sample2[9] ),
    .A2(_03424_),
    .B(_07565_),
    .C(_03233_),
    .ZN(_07566_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15634_ (.A1(\channels.sample1[9] ),
    .A2(_03427_),
    .ZN(_07567_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _15635_ (.A1(_07566_),
    .A2(_07567_),
    .ZN(_07568_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _15636_ (.A1(\filters.sample_buff[9] ),
    .A2(_07568_),
    .Z(_07569_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _15637_ (.A1(_07562_),
    .A2(_07557_),
    .A3(_07569_),
    .Z(_07570_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _15638_ (.A1(_07562_),
    .A2(_07557_),
    .B(_07569_),
    .ZN(_07571_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15639_ (.A1(_07486_),
    .A2(_07570_),
    .A3(_07571_),
    .ZN(_07572_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15640_ (.I(_06978_),
    .Z(_07573_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15641_ (.A1(_07561_),
    .A2(_07572_),
    .B(_07573_),
    .ZN(_00599_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15642_ (.A1(\filters.sample_buff[9] ),
    .A2(_07568_),
    .ZN(_07574_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15643_ (.A1(\channels.sample3[10] ),
    .A2(_07549_),
    .ZN(_07575_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _15644_ (.A1(_03409_),
    .A2(_07563_),
    .B(_07575_),
    .C(_03424_),
    .ZN(_07576_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _15645_ (.A1(\channels.sample2[10] ),
    .A2(_03424_),
    .B(_07576_),
    .C(_03234_),
    .ZN(_07577_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15646_ (.A1(\channels.sample1[10] ),
    .A2(_03428_),
    .ZN(_07578_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15647_ (.A1(_07577_),
    .A2(_07578_),
    .ZN(_07579_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _15648_ (.A1(\filters.sample_buff[10] ),
    .A2(_07579_),
    .Z(_07580_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _15649_ (.I(_07580_),
    .ZN(_07581_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _15650_ (.A1(_07574_),
    .A2(_07571_),
    .B(_07581_),
    .ZN(_07582_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _15651_ (.A1(_07574_),
    .A2(_07571_),
    .A3(_07581_),
    .Z(_07583_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15652_ (.A1(_07582_),
    .A2(_07583_),
    .ZN(_07584_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _15653_ (.A1(\filters.sample_buff[10] ),
    .A2(_07447_),
    .B1(_07523_),
    .B2(_07584_),
    .ZN(_07585_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15654_ (.A1(_07498_),
    .A2(_07585_),
    .ZN(_00600_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15655_ (.A1(\filters.sample_buff[11] ),
    .A2(_07448_),
    .ZN(_07586_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _15656_ (.A1(\filters.sample_buff[10] ),
    .A2(_07579_),
    .Z(_07587_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15657_ (.A1(_02056_),
    .A2(_07563_),
    .ZN(_07588_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _15658_ (.A1(_03421_),
    .A2(_07563_),
    .B(_07588_),
    .C(_03224_),
    .ZN(_07589_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _15659_ (.A1(\channels.sample2[11] ),
    .A2(_03225_),
    .B(_07589_),
    .C(_03234_),
    .ZN(_07590_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15660_ (.A1(\channels.sample1[11] ),
    .A2(_03428_),
    .ZN(_07591_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15661_ (.A1(_07590_),
    .A2(_07591_),
    .ZN(_07592_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _15662_ (.A1(\filters.sample_buff[11] ),
    .A2(_07592_),
    .Z(_07593_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _15663_ (.A1(_07587_),
    .A2(_07582_),
    .A3(_07593_),
    .Z(_07594_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15664_ (.A1(_07587_),
    .A2(_07582_),
    .B(_07593_),
    .ZN(_07595_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15665_ (.A1(_07450_),
    .A2(_07594_),
    .A3(_07595_),
    .ZN(_07596_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15666_ (.A1(_07586_),
    .A2(_07596_),
    .B(_07573_),
    .ZN(_00601_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _15667_ (.I(_03940_),
    .Z(_07597_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _15668_ (.I(_07597_),
    .Z(_07598_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15669_ (.A1(\filters.sample_buff[11] ),
    .A2(_07592_),
    .ZN(_07599_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15670_ (.A1(_07599_),
    .A2(_07595_),
    .ZN(_07600_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15671_ (.A1(_03239_),
    .A2(_03237_),
    .ZN(_07601_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _15672_ (.I(_07601_),
    .Z(_07602_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _15673_ (.A1(\filters.sample_buff[12] ),
    .A2(_03450_),
    .A3(_07602_),
    .Z(_07603_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15674_ (.A1(_03450_),
    .A2(_07602_),
    .B(\filters.sample_buff[12] ),
    .ZN(_07604_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15675_ (.A1(_07603_),
    .A2(_07604_),
    .ZN(_07605_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _15676_ (.A1(_07600_),
    .A2(_07605_),
    .Z(_07606_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _15677_ (.A1(\filters.sample_buff[12] ),
    .A2(_07447_),
    .B1(_07523_),
    .B2(_07606_),
    .ZN(_07607_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15678_ (.A1(_07598_),
    .A2(_07607_),
    .ZN(_00602_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15679_ (.A1(\filters.sample_buff[13] ),
    .A2(_07448_),
    .ZN(_07608_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _15680_ (.A1(_07600_),
    .A2(_07605_),
    .Z(_07609_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15681_ (.A1(\filters.sample_filtered[14] ),
    .A2(_07601_),
    .ZN(_07610_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _15682_ (.A1(\filters.sample_buff[13] ),
    .A2(_07610_),
    .ZN(_07611_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _15683_ (.A1(_07603_),
    .A2(_07609_),
    .A3(_07611_),
    .Z(_07612_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _15684_ (.A1(_07603_),
    .A2(_07609_),
    .B(_07611_),
    .ZN(_07613_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15685_ (.A1(_07450_),
    .A2(_07612_),
    .A3(_07613_),
    .ZN(_07614_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15686_ (.A1(_07608_),
    .A2(_07614_),
    .B(_07573_),
    .ZN(_00603_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _15687_ (.I(\filters.sample_buff[14] ),
    .ZN(_07615_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15688_ (.A1(\filters.sample_buff[13] ),
    .A2(_03452_),
    .A3(_07602_),
    .ZN(_07616_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15689_ (.A1(\filters.sample_filtered[15] ),
    .A2(_07602_),
    .ZN(_07617_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _15690_ (.A1(_07615_),
    .A2(_07617_),
    .Z(_07618_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15691_ (.A1(_07616_),
    .A2(_07613_),
    .B(_07618_),
    .ZN(_07619_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15692_ (.A1(_07616_),
    .A2(_07613_),
    .A3(_07618_),
    .ZN(_07620_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15693_ (.A1(_07450_),
    .A2(_07620_),
    .ZN(_07621_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15694_ (.A1(_07619_),
    .A2(_07621_),
    .ZN(_07622_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _15695_ (.A1(_07615_),
    .A2(_07484_),
    .B(_07622_),
    .C(_07269_),
    .ZN(_00604_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _15696_ (.I(\channels.exp_periods[3][0] ),
    .Z(_07623_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _15697_ (.I(_07623_),
    .Z(_00605_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _15698_ (.I(\channels.exp_periods[3][1] ),
    .Z(_07624_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _15699_ (.I(_07624_),
    .Z(_00606_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _15700_ (.I(\channels.exp_periods[3][2] ),
    .Z(_07625_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _15701_ (.I(_07625_),
    .Z(_00607_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _15702_ (.I(\channels.exp_periods[3][3] ),
    .Z(_07626_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _15703_ (.I(_07626_),
    .Z(_00608_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _15704_ (.I(\channels.exp_periods[3][4] ),
    .Z(_07627_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _15705_ (.I(_07627_),
    .Z(_00609_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15706_ (.A1(_03216_),
    .A2(_03729_),
    .ZN(_07628_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _15707_ (.A1(_07443_),
    .A2(_03214_),
    .A3(_07628_),
    .ZN(_07629_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _15708_ (.I(_07629_),
    .Z(_07630_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _15709_ (.I(_07630_),
    .Z(_07631_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _15710_ (.I(_07631_),
    .Z(_07632_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15711_ (.I(_07630_),
    .Z(_07633_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15712_ (.A1(_05534_),
    .A2(_07633_),
    .B(_07356_),
    .ZN(_07634_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15713_ (.A1(_05539_),
    .A2(_07632_),
    .B(_07634_),
    .ZN(_00610_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15714_ (.A1(_03216_),
    .A2(_03730_),
    .A3(_03205_),
    .ZN(_07635_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _15715_ (.I(_07635_),
    .Z(_07636_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15716_ (.I(_07636_),
    .Z(_07637_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15717_ (.A1(_05651_),
    .A2(_07637_),
    .ZN(_07638_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _15718_ (.I(_07629_),
    .Z(_07639_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _15719_ (.I(_07639_),
    .Z(_07640_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15720_ (.A1(_05647_),
    .A2(_07640_),
    .B(_07333_),
    .ZN(_07641_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15721_ (.A1(_07638_),
    .A2(_07641_),
    .ZN(_00611_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15722_ (.A1(_05759_),
    .A2(_07637_),
    .ZN(_07642_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15723_ (.I(_07639_),
    .Z(_07643_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15724_ (.I(_07332_),
    .Z(_07644_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15725_ (.A1(_03268_),
    .A2(_07643_),
    .B(_07644_),
    .ZN(_07645_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15726_ (.A1(_07642_),
    .A2(_07645_),
    .ZN(_00612_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15727_ (.A1(_05862_),
    .A2(_07637_),
    .ZN(_07646_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15728_ (.A1(_03282_),
    .A2(_07643_),
    .B(_07644_),
    .ZN(_07647_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15729_ (.A1(_07646_),
    .A2(_07647_),
    .ZN(_00613_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _15730_ (.I(_07355_),
    .Z(_07648_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15731_ (.A1(_05969_),
    .A2(_07633_),
    .B(_07648_),
    .ZN(_07649_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15732_ (.A1(_05973_),
    .A2(_07632_),
    .B(_07649_),
    .ZN(_00614_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15733_ (.A1(_06078_),
    .A2(_07637_),
    .ZN(_07650_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15734_ (.A1(_03310_),
    .A2(_07643_),
    .B(_07644_),
    .ZN(_07651_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15735_ (.A1(_07650_),
    .A2(_07651_),
    .ZN(_00615_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15736_ (.I(_07636_),
    .Z(_07652_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15737_ (.A1(_06184_),
    .A2(_07652_),
    .ZN(_07653_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15738_ (.A1(_03329_),
    .A2(_07643_),
    .B(_07644_),
    .ZN(_07654_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15739_ (.A1(_07653_),
    .A2(_07654_),
    .ZN(_00616_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15740_ (.A1(_06291_),
    .A2(_07652_),
    .ZN(_07655_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15741_ (.I(_07639_),
    .Z(_07656_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15742_ (.I(_07332_),
    .Z(_07657_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15743_ (.A1(_03345_),
    .A2(_07656_),
    .B(_07657_),
    .ZN(_07658_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15744_ (.A1(_07655_),
    .A2(_07658_),
    .ZN(_00617_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15745_ (.A1(_06401_),
    .A2(_07652_),
    .ZN(_07659_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15746_ (.A1(_03360_),
    .A2(_07656_),
    .B(_07657_),
    .ZN(_07660_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15747_ (.A1(_07659_),
    .A2(_07660_),
    .ZN(_00618_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15748_ (.A1(_06506_),
    .A2(_07652_),
    .ZN(_07661_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15749_ (.A1(_03374_),
    .A2(_07656_),
    .B(_07657_),
    .ZN(_07662_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15750_ (.A1(_07661_),
    .A2(_07662_),
    .ZN(_00619_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _15751_ (.I(_07635_),
    .Z(_07663_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15752_ (.I(_07663_),
    .Z(_07664_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15753_ (.A1(_06608_),
    .A2(_07664_),
    .ZN(_07665_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15754_ (.A1(_03394_),
    .A2(_07656_),
    .B(_07657_),
    .ZN(_07666_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15755_ (.A1(_07665_),
    .A2(_07666_),
    .ZN(_00620_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15756_ (.A1(_03411_),
    .A2(_07633_),
    .B(_07648_),
    .ZN(_07667_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15757_ (.A1(_06695_),
    .A2(_07632_),
    .B(_07667_),
    .ZN(_00621_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15758_ (.A1(_03422_),
    .A2(_07633_),
    .B(_07648_),
    .ZN(_07668_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15759_ (.A1(_06714_),
    .A2(_07632_),
    .B(_07668_),
    .ZN(_00622_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15760_ (.A1(_06728_),
    .A2(_07664_),
    .ZN(_07669_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _15761_ (.I(_07639_),
    .Z(_07670_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _15762_ (.I(_07332_),
    .Z(_07671_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15763_ (.A1(_03439_),
    .A2(_07670_),
    .B(_07671_),
    .ZN(_07672_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15764_ (.A1(_07669_),
    .A2(_07672_),
    .ZN(_00623_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15765_ (.A1(_06737_),
    .A2(_07664_),
    .ZN(_07673_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15766_ (.A1(_03455_),
    .A2(_07670_),
    .B(_07671_),
    .ZN(_07674_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15767_ (.A1(_07673_),
    .A2(_07674_),
    .ZN(_00624_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15768_ (.A1(_06746_),
    .A2(_07664_),
    .ZN(_07675_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15769_ (.A1(_03468_),
    .A2(_07670_),
    .B(_07671_),
    .ZN(_07676_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15770_ (.A1(_07675_),
    .A2(_07676_),
    .ZN(_00625_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15771_ (.I(_07663_),
    .Z(_07677_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15772_ (.A1(_06758_),
    .A2(_07677_),
    .ZN(_07678_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15773_ (.A1(\filters.low[16] ),
    .A2(_07670_),
    .B(_07671_),
    .ZN(_07679_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15774_ (.A1(_07678_),
    .A2(_07679_),
    .ZN(_00626_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15775_ (.A1(_07295_),
    .A2(_07631_),
    .B(_07648_),
    .ZN(_07680_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15776_ (.A1(_06774_),
    .A2(_07640_),
    .B(_07680_),
    .ZN(_00627_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15777_ (.A1(_06783_),
    .A2(_07677_),
    .ZN(_07681_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15778_ (.I(_07630_),
    .Z(_07682_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _15779_ (.I(_03733_),
    .Z(_07683_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _15780_ (.I(_07683_),
    .Z(_07684_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15781_ (.A1(\filters.low[18] ),
    .A2(_07682_),
    .B(_07684_),
    .ZN(_07685_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15782_ (.A1(_07681_),
    .A2(_07685_),
    .ZN(_00628_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15783_ (.A1(_06791_),
    .A2(_07677_),
    .ZN(_07686_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15784_ (.A1(\filters.low[19] ),
    .A2(_07682_),
    .B(_07684_),
    .ZN(_07687_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15785_ (.A1(_07686_),
    .A2(_07687_),
    .ZN(_00629_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15786_ (.A1(_06801_),
    .A2(_07677_),
    .ZN(_07688_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15787_ (.A1(\filters.low[20] ),
    .A2(_07682_),
    .B(_07684_),
    .ZN(_07689_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15788_ (.A1(_07688_),
    .A2(_07689_),
    .ZN(_00630_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15789_ (.I(_07663_),
    .Z(_07690_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15790_ (.A1(_06809_),
    .A2(_07690_),
    .ZN(_07691_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15791_ (.A1(_07327_),
    .A2(_07682_),
    .B(_07684_),
    .ZN(_07692_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15792_ (.A1(_07691_),
    .A2(_07692_),
    .ZN(_00631_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15793_ (.A1(_06818_),
    .A2(_07690_),
    .ZN(_07693_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15794_ (.I(_07630_),
    .Z(_07694_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15795_ (.I(_07683_),
    .Z(_07695_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15796_ (.A1(\filters.low[22] ),
    .A2(_07694_),
    .B(_07695_),
    .ZN(_07696_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15797_ (.A1(_07693_),
    .A2(_07696_),
    .ZN(_00632_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15798_ (.I(_07636_),
    .Z(_07697_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15799_ (.I(_07663_),
    .Z(_07698_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15800_ (.A1(_06828_),
    .A2(_07698_),
    .ZN(_07699_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _15801_ (.A1(_06822_),
    .A2(_07697_),
    .B(_07699_),
    .C(_07269_),
    .ZN(_00633_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _15802_ (.I(_07355_),
    .Z(_07700_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15803_ (.A1(_07363_),
    .A2(_07631_),
    .B(_07700_),
    .ZN(_07701_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15804_ (.A1(_06841_),
    .A2(_07640_),
    .B(_07701_),
    .ZN(_00634_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15805_ (.A1(_06848_),
    .A2(_07690_),
    .ZN(_07702_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15806_ (.A1(_07373_),
    .A2(_07694_),
    .B(_07695_),
    .ZN(_07703_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15807_ (.A1(_07702_),
    .A2(_07703_),
    .ZN(_00635_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15808_ (.A1(_06858_),
    .A2(_07690_),
    .ZN(_07704_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15809_ (.A1(_07383_),
    .A2(_07694_),
    .B(_07695_),
    .ZN(_07705_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15810_ (.A1(_07704_),
    .A2(_07705_),
    .ZN(_00636_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15811_ (.A1(_06867_),
    .A2(_07698_),
    .ZN(_07706_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15812_ (.A1(_07395_),
    .A2(_07694_),
    .B(_07695_),
    .ZN(_07707_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15813_ (.A1(_07706_),
    .A2(_07707_),
    .ZN(_00637_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15814_ (.A1(_06879_),
    .A2(_07698_),
    .ZN(_07708_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _15815_ (.A1(_06875_),
    .A2(_07697_),
    .B(_07708_),
    .C(_07269_),
    .ZN(_00638_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15816_ (.A1(_06888_),
    .A2(_07698_),
    .ZN(_07709_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _15817_ (.I(_02353_),
    .Z(_07710_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _15818_ (.A1(_06882_),
    .A2(_07697_),
    .B(_07709_),
    .C(_07710_),
    .ZN(_00639_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15819_ (.A1(_06897_),
    .A2(_07636_),
    .ZN(_07711_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _15820_ (.A1(_06891_),
    .A2(_07697_),
    .B(_07711_),
    .C(_07710_),
    .ZN(_00640_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15821_ (.A1(\filters.low[31] ),
    .A2(_07631_),
    .B(_07700_),
    .ZN(_07712_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15822_ (.A1(_06905_),
    .A2(_07640_),
    .B(_07712_),
    .ZN(_00641_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15823_ (.A1(_03735_),
    .A2(_07628_),
    .ZN(_07713_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _15824_ (.A1(_04189_),
    .A2(_04158_),
    .B(_07713_),
    .ZN(_00642_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15825_ (.A1(_03214_),
    .A2(_03216_),
    .A3(_03731_),
    .ZN(_07714_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15826_ (.A1(_03735_),
    .A2(_07714_),
    .ZN(_07715_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _15827_ (.A1(_03194_),
    .A2(_07628_),
    .B(_07715_),
    .ZN(_00643_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _15828_ (.A1(_07443_),
    .A2(_07714_),
    .Z(_07716_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _15829_ (.A1(_07598_),
    .A2(_07716_),
    .ZN(_00644_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _15830_ (.A1(\spi_dac_i.counter[4] ),
    .A2(\spi_dac_i.counter[3] ),
    .Z(_07717_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _15831_ (.A1(\spi_dac_i.counter[0] ),
    .A2(_07717_),
    .Z(_07718_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15832_ (.I(_07718_),
    .Z(_07719_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15833_ (.I(\spi_dac_i.counter[0] ),
    .Z(_07720_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15834_ (.I(_07717_),
    .Z(_07721_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _15835_ (.I(_07721_),
    .Z(_07722_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15836_ (.A1(_07720_),
    .A2(_04776_),
    .A3(_07722_),
    .ZN(_07723_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15837_ (.A1(_07719_),
    .A2(_07723_),
    .B(_07573_),
    .ZN(_00645_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15838_ (.I(\spi_dac_i.counter[3] ),
    .Z(_07724_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15839_ (.A1(\spi_dac_i.counter[4] ),
    .A2(_07724_),
    .ZN(_07725_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15840_ (.I(_07725_),
    .Z(_07726_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _15841_ (.A1(\spi_dac_i.counter[0] ),
    .A2(_07726_),
    .Z(_07727_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _15842_ (.I(_07727_),
    .Z(_07728_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _15843_ (.I(_07718_),
    .Z(_07729_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15844_ (.A1(_04776_),
    .A2(_07721_),
    .ZN(_07730_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15845_ (.A1(\spi_dac_i.counter[1] ),
    .A2(_07729_),
    .A3(_07730_),
    .ZN(_07731_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15846_ (.A1(\spi_dac_i.counter[1] ),
    .A2(_07728_),
    .B(_07731_),
    .ZN(_07732_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15847_ (.A1(_07598_),
    .A2(_07732_),
    .ZN(_00646_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _15848_ (.A1(\spi_dac_i.counter[2] ),
    .A2(\spi_dac_i.counter[1] ),
    .A3(_07720_),
    .Z(_07733_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15849_ (.A1(\spi_dac_i.counter[1] ),
    .A2(_07720_),
    .B(\spi_dac_i.counter[2] ),
    .ZN(_07734_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _15850_ (.I(\spi_dac_i.counter[2] ),
    .ZN(_07735_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _15851_ (.A1(_07721_),
    .A2(_07733_),
    .A3(_07734_),
    .B1(_07730_),
    .B2(_07735_),
    .ZN(_07736_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _15852_ (.A1(_03735_),
    .A2(_07736_),
    .Z(_07737_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _15853_ (.I(_07737_),
    .Z(_00647_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15854_ (.A1(\spi_dac_i.counter[4] ),
    .A2(_07733_),
    .B(_07724_),
    .ZN(_07738_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15855_ (.A1(_07724_),
    .A2(_07733_),
    .B(_07738_),
    .ZN(_07739_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _15856_ (.I(_01822_),
    .Z(_07740_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15857_ (.A1(_07730_),
    .A2(_07739_),
    .B(_07740_),
    .ZN(_00648_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15858_ (.I(_07717_),
    .Z(_07741_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _15859_ (.I(_07741_),
    .Z(_07742_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15860_ (.I(_07742_),
    .Z(_07743_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15861_ (.A1(_07724_),
    .A2(_07733_),
    .B(\spi_dac_i.counter[4] ),
    .ZN(_07744_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _15862_ (.A1(_04170_),
    .A2(_07743_),
    .B(_07744_),
    .C(_07710_),
    .ZN(_00649_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _15863_ (.I(\tt_um_rejunity_sn76489.chan[2].attenuation.in ),
    .ZN(_07745_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _15864_ (.I(_07745_),
    .Z(_07746_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _15865_ (.A1(\tt_um_rejunity_sn76489.chan[2].attenuation.control[3] ),
    .A2(_07746_),
    .ZN(_07747_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _15866_ (.A1(\tt_um_rejunity_sn76489.chan[2].attenuation.control[2] ),
    .A2(_07746_),
    .ZN(_07748_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15867_ (.I(_07748_),
    .Z(_07749_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15868_ (.A1(\tt_um_rejunity_sn76489.chan[2].attenuation.control[1] ),
    .A2(_07745_),
    .ZN(_07750_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _15869_ (.I(_07750_),
    .Z(_07751_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15870_ (.A1(\tt_um_rejunity_sn76489.chan[2].attenuation.control[0] ),
    .A2(_07749_),
    .ZN(_07752_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _15871_ (.A1(_07749_),
    .A2(_07751_),
    .B(_07752_),
    .ZN(_07753_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _15872_ (.A1(\tt_um_rejunity_sn76489.chan[2].attenuation.control[0] ),
    .A2(_07746_),
    .ZN(_07754_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _15873_ (.I(\tt_um_rejunity_sn76489.chan[2].attenuation.control[2] ),
    .ZN(_07755_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15874_ (.A1(_07755_),
    .A2(\tt_um_rejunity_sn76489.chan[2].attenuation.in ),
    .ZN(_07756_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15875_ (.I(_07756_),
    .Z(_07757_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _15876_ (.A1(_07757_),
    .A2(_07751_),
    .Z(_07758_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _15877_ (.I(\tt_um_rejunity_sn76489.chan[2].attenuation.control[3] ),
    .ZN(_07759_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _15878_ (.A1(_07759_),
    .A2(_02347_),
    .ZN(_07760_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15879_ (.I(_07760_),
    .Z(_07761_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15880_ (.A1(_07754_),
    .A2(_07758_),
    .B(_07761_),
    .ZN(_07762_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _15881_ (.I(_07762_),
    .ZN(_07763_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15882_ (.A1(_07747_),
    .A2(_07753_),
    .B(_07763_),
    .ZN(_07764_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _15883_ (.I(\tt_um_rejunity_sn76489.chan[1].attenuation.in ),
    .ZN(_07765_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15884_ (.I(_07765_),
    .Z(_07766_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _15885_ (.A1(\tt_um_rejunity_sn76489.chan[1].attenuation.control[3] ),
    .A2(_07766_),
    .ZN(_07767_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15886_ (.A1(\tt_um_rejunity_sn76489.chan[1].attenuation.control[2] ),
    .A2(_07765_),
    .ZN(_07768_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _15887_ (.A1(\tt_um_rejunity_sn76489.chan[1].attenuation.control[1] ),
    .A2(_07766_),
    .ZN(_07769_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15888_ (.A1(\tt_um_rejunity_sn76489.chan[1].attenuation.control[0] ),
    .A2(_07768_),
    .ZN(_07770_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15889_ (.A1(_07768_),
    .A2(_07769_),
    .B(_07770_),
    .ZN(_07771_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _15890_ (.A1(\tt_um_rejunity_sn76489.chan[1].attenuation.control[2] ),
    .A2(_07765_),
    .Z(_07772_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15891_ (.I(_07772_),
    .Z(_07773_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _15892_ (.I(\tt_um_rejunity_sn76489.chan[1].attenuation.control[1] ),
    .ZN(_07774_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15893_ (.A1(_07774_),
    .A2(\tt_um_rejunity_sn76489.chan[1].attenuation.in ),
    .ZN(_07775_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _15894_ (.A1(_07773_),
    .A2(_07775_),
    .ZN(_07776_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _15895_ (.I(_07768_),
    .Z(_07777_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _15896_ (.A1(\tt_um_rejunity_sn76489.chan[1].attenuation.control[0] ),
    .A2(_07766_),
    .Z(_07778_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15897_ (.A1(_07777_),
    .A2(_07769_),
    .B(_07778_),
    .ZN(_07779_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _15898_ (.A1(\tt_um_rejunity_sn76489.chan[1].attenuation.control[3] ),
    .A2(_07766_),
    .Z(_07780_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _15899_ (.A1(_07776_),
    .A2(_07779_),
    .B(_07780_),
    .ZN(_07781_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _15900_ (.I(_07781_),
    .ZN(_07782_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15901_ (.A1(_07767_),
    .A2(_07771_),
    .B(_07782_),
    .ZN(_07783_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _15902_ (.I(\tt_um_rejunity_sn76489.chan[0].attenuation.control[2] ),
    .ZN(_07784_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15903_ (.A1(_07784_),
    .A2(\tt_um_rejunity_sn76489.chan[0].attenuation.in ),
    .ZN(_07785_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15904_ (.I(_07785_),
    .Z(_07786_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _15905_ (.I(\tt_um_rejunity_sn76489.chan[0].attenuation.in ),
    .ZN(_07787_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _15906_ (.A1(\tt_um_rejunity_sn76489.chan[0].attenuation.control[1] ),
    .A2(_07787_),
    .ZN(_07788_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15907_ (.A1(_07786_),
    .A2(_07788_),
    .ZN(_07789_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15908_ (.I(_07787_),
    .Z(_07790_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15909_ (.A1(\tt_um_rejunity_sn76489.chan[0].attenuation.control[2] ),
    .A2(_07790_),
    .ZN(_07791_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _15910_ (.I(_07791_),
    .Z(_07792_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15911_ (.A1(\tt_um_rejunity_sn76489.chan[0].attenuation.control[0] ),
    .A2(_07790_),
    .ZN(_07793_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15912_ (.I(_07793_),
    .Z(_07794_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _15913_ (.A1(\tt_um_rejunity_sn76489.chan[0].attenuation.control[3] ),
    .A2(_07790_),
    .Z(_07795_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15914_ (.A1(_07792_),
    .A2(_07794_),
    .B(_07795_),
    .ZN(_07796_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _15915_ (.I(\tt_um_rejunity_sn76489.chan[0].attenuation.control[1] ),
    .ZN(_07797_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15916_ (.I(\tt_um_rejunity_sn76489.chan[0].attenuation.in ),
    .Z(_07798_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15917_ (.A1(_07797_),
    .A2(_07798_),
    .ZN(_07799_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _15918_ (.A1(_07785_),
    .A2(_07799_),
    .ZN(_07800_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15919_ (.I(\tt_um_rejunity_sn76489.chan[0].attenuation.control[0] ),
    .Z(_07801_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _15920_ (.A1(_07784_),
    .A2(_07797_),
    .B(_07801_),
    .C(_07798_),
    .ZN(_07802_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15921_ (.A1(_07800_),
    .A2(_07802_),
    .B(_07795_),
    .ZN(_07803_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _15922_ (.I(_07803_),
    .ZN(_07804_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15923_ (.A1(_07789_),
    .A2(_07796_),
    .B(_07804_),
    .ZN(_07805_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _15924_ (.A1(_07783_),
    .A2(_07805_),
    .ZN(_07806_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _15925_ (.I(_07806_),
    .ZN(_07807_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _15926_ (.I(\tt_um_rejunity_sn76489.chan[3].attenuation.in ),
    .ZN(_07808_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15927_ (.I(_07808_),
    .Z(_07809_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _15928_ (.A1(\tt_um_rejunity_sn76489.chan[3].attenuation.control[3] ),
    .A2(_07809_),
    .ZN(_07810_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _15929_ (.I(_07810_),
    .Z(_07811_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15930_ (.A1(\tt_um_rejunity_sn76489.chan[3].attenuation.control[2] ),
    .A2(_07808_),
    .ZN(_07812_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15931_ (.I(_07812_),
    .Z(_07813_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _15932_ (.A1(\tt_um_rejunity_sn76489.chan[3].attenuation.control[1] ),
    .A2(_07809_),
    .ZN(_07814_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15933_ (.A1(\tt_um_rejunity_sn76489.chan[3].attenuation.control[0] ),
    .A2(_07812_),
    .ZN(_07815_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _15934_ (.A1(_07813_),
    .A2(_07814_),
    .B(_07815_),
    .ZN(_07816_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _15935_ (.I(\tt_um_rejunity_sn76489.chan[3].attenuation.control[2] ),
    .ZN(_07817_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _15936_ (.I(\tt_um_rejunity_sn76489.chan[3].attenuation.in ),
    .Z(_07818_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15937_ (.A1(_07817_),
    .A2(_07818_),
    .ZN(_07819_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15938_ (.I(_07819_),
    .Z(_07820_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _15939_ (.I(\tt_um_rejunity_sn76489.chan[3].attenuation.control[1] ),
    .ZN(_07821_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15940_ (.A1(_07821_),
    .A2(_07818_),
    .ZN(_07822_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _15941_ (.I(_07822_),
    .Z(_07823_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15942_ (.A1(_07820_),
    .A2(_07823_),
    .ZN(_07824_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _15943_ (.I(_07813_),
    .Z(_07825_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _15944_ (.I(\tt_um_rejunity_sn76489.chan[3].attenuation.control[0] ),
    .ZN(_07826_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _15945_ (.A1(_07826_),
    .A2(\tt_um_rejunity_sn76489.chan[3].attenuation.in ),
    .ZN(_07827_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15946_ (.A1(_07825_),
    .A2(_07814_),
    .B(_07827_),
    .ZN(_07828_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15947_ (.A1(_07824_),
    .A2(_07828_),
    .ZN(_07829_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15948_ (.A1(_07810_),
    .A2(_07829_),
    .ZN(_07830_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _15949_ (.A1(_07811_),
    .A2(_07816_),
    .B(_07830_),
    .ZN(_07831_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _15950_ (.A1(_07807_),
    .A2(_07831_),
    .Z(_07832_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15951_ (.A1(_07764_),
    .A2(_07832_),
    .ZN(_07833_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15952_ (.I(_07726_),
    .Z(_07834_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15953_ (.A1(_07764_),
    .A2(_07832_),
    .ZN(_07835_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15954_ (.A1(_07834_),
    .A2(_07835_),
    .ZN(_07836_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _15955_ (.A1(\spi_dac_i.spi_dat_buff_1[0] ),
    .A2(_07728_),
    .B1(_07833_),
    .B2(_07836_),
    .ZN(_07837_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15956_ (.A1(_07598_),
    .A2(_07837_),
    .ZN(_00650_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _15957_ (.I(_07722_),
    .Z(_07838_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15958_ (.A1(_07807_),
    .A2(_07831_),
    .ZN(_07839_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15959_ (.A1(_07839_),
    .A2(_07833_),
    .ZN(_07840_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _15960_ (.I(\tt_um_rejunity_sn76489.chan[2].attenuation.control[1] ),
    .Z(_07841_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15961_ (.A1(_07747_),
    .A2(_07752_),
    .ZN(_07842_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15962_ (.A1(_07757_),
    .A2(_07754_),
    .ZN(_07843_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15963_ (.A1(_07761_),
    .A2(_07843_),
    .ZN(_07844_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _15964_ (.A1(_07841_),
    .A2(_07842_),
    .B1(_07844_),
    .B2(_07753_),
    .ZN(_07845_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15965_ (.A1(_07813_),
    .A2(_07827_),
    .ZN(_07846_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15966_ (.A1(_07810_),
    .A2(_07815_),
    .ZN(_07847_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _15967_ (.A1(_07810_),
    .A2(_07816_),
    .A3(_07846_),
    .B1(_07847_),
    .B2(\tt_um_rejunity_sn76489.chan[3].attenuation.control[1] ),
    .ZN(_07848_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _15968_ (.A1(_07783_),
    .A2(_07805_),
    .Z(_07849_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15969_ (.A1(_07801_),
    .A2(_07791_),
    .ZN(_07850_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15970_ (.A1(\tt_um_rejunity_sn76489.chan[0].attenuation.control[0] ),
    .A2(_07788_),
    .ZN(_07851_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15971_ (.A1(_07795_),
    .A2(_07786_),
    .A3(_07851_),
    .ZN(_07852_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _15972_ (.A1(\tt_um_rejunity_sn76489.chan[0].attenuation.control[3] ),
    .A2(_07790_),
    .ZN(_07853_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15973_ (.A1(\tt_um_rejunity_sn76489.chan[0].attenuation.control[1] ),
    .A2(_07853_),
    .ZN(_07854_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15974_ (.A1(_07850_),
    .A2(_07852_),
    .A3(_07854_),
    .ZN(_07855_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15975_ (.A1(_07767_),
    .A2(_07770_),
    .ZN(_07856_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15976_ (.A1(\tt_um_rejunity_sn76489.chan[1].attenuation.control[0] ),
    .A2(_07765_),
    .ZN(_07857_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15977_ (.A1(_07772_),
    .A2(_07857_),
    .ZN(_07858_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15978_ (.A1(_07780_),
    .A2(_07858_),
    .ZN(_07859_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _15979_ (.A1(\tt_um_rejunity_sn76489.chan[1].attenuation.control[1] ),
    .A2(_07856_),
    .B1(_07859_),
    .B2(_07771_),
    .ZN(_07860_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _15980_ (.A1(_07855_),
    .A2(_07860_),
    .Z(_07861_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _15981_ (.I(_07861_),
    .ZN(_07862_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _15982_ (.A1(_07849_),
    .A2(_07862_),
    .Z(_07863_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _15983_ (.A1(_07848_),
    .A2(_07863_),
    .Z(_07864_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _15984_ (.A1(_07845_),
    .A2(_07864_),
    .ZN(_07865_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _15985_ (.A1(_07840_),
    .A2(_07865_),
    .Z(_07866_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15986_ (.I(_07729_),
    .Z(_07867_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15987_ (.A1(\spi_dac_i.counter[0] ),
    .A2(_07725_),
    .ZN(_07868_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _15988_ (.I(_07868_),
    .Z(_07869_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15989_ (.I(_07869_),
    .Z(_07870_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15990_ (.I(_02101_),
    .Z(_07871_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _15991_ (.A1(\spi_dac_i.spi_dat_buff_1[0] ),
    .A2(_07867_),
    .B1(_07870_),
    .B2(\spi_dac_i.spi_dat_buff_1[1] ),
    .C(_07871_),
    .ZN(_07872_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15992_ (.A1(_07838_),
    .A2(_07866_),
    .B(_07872_),
    .ZN(_00651_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15993_ (.A1(_07839_),
    .A2(_07833_),
    .B(_07865_),
    .ZN(_07873_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _15994_ (.A1(_07750_),
    .A2(_07754_),
    .ZN(_07874_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _15995_ (.I(_07874_),
    .Z(_07875_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _15996_ (.A1(_07841_),
    .A2(\tt_um_rejunity_sn76489.chan[2].attenuation.control[0] ),
    .A3(_07746_),
    .ZN(_07876_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _15997_ (.A1(_07748_),
    .A2(_07874_),
    .A3(_07876_),
    .ZN(_07877_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _15998_ (.A1(_07756_),
    .A2(_07751_),
    .ZN(_07878_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _15999_ (.A1(_07747_),
    .A2(_07878_),
    .ZN(_07879_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _16000_ (.A1(_07748_),
    .A2(_07875_),
    .B(_07877_),
    .C(_07879_),
    .ZN(_07880_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _16001_ (.A1(_07788_),
    .A2(_07794_),
    .ZN(_07881_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _16002_ (.A1(_07788_),
    .A2(_07793_),
    .ZN(_07882_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16003_ (.A1(_07792_),
    .A2(_07882_),
    .ZN(_07883_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16004_ (.A1(_07881_),
    .A2(_07883_),
    .ZN(_07884_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16005_ (.A1(_07799_),
    .A2(_07794_),
    .ZN(_07885_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16006_ (.A1(_07791_),
    .A2(_07799_),
    .ZN(_07886_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _16007_ (.A1(_07853_),
    .A2(_07886_),
    .ZN(_07887_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16008_ (.A1(_07885_),
    .A2(_07887_),
    .ZN(_07888_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16009_ (.A1(_07884_),
    .A2(_07888_),
    .ZN(_07889_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _16010_ (.I(_07775_),
    .Z(_07890_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16011_ (.A1(_07890_),
    .A2(_07778_),
    .ZN(_07891_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _16012_ (.A1(_07769_),
    .A2(_07857_),
    .Z(_07892_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _16013_ (.A1(_07777_),
    .A2(_07890_),
    .B(_07767_),
    .ZN(_07893_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16014_ (.A1(_07773_),
    .A2(_07892_),
    .B(_07893_),
    .ZN(_07894_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16015_ (.A1(_07773_),
    .A2(_07891_),
    .B(_07894_),
    .ZN(_07895_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16016_ (.A1(_07889_),
    .A2(_07895_),
    .ZN(_07896_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _16017_ (.I(_07896_),
    .ZN(_07897_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16018_ (.A1(_07889_),
    .A2(_07895_),
    .ZN(_07898_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16019_ (.A1(_07897_),
    .A2(_07898_),
    .ZN(_07899_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _16020_ (.A1(_07850_),
    .A2(_07852_),
    .A3(_07854_),
    .A4(_07860_),
    .ZN(_07900_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16021_ (.A1(_07849_),
    .A2(_07862_),
    .ZN(_07901_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _16022_ (.A1(_07900_),
    .A2(_07901_),
    .ZN(_07902_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _16023_ (.A1(_07899_),
    .A2(_07902_),
    .ZN(_07903_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16024_ (.A1(_07822_),
    .A2(_07827_),
    .ZN(_07904_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16025_ (.A1(\tt_um_rejunity_sn76489.chan[3].attenuation.control[0] ),
    .A2(_07809_),
    .ZN(_07905_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16026_ (.A1(_07814_),
    .A2(_07905_),
    .ZN(_07906_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _16027_ (.A1(_07904_),
    .A2(_07906_),
    .Z(_07907_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _16028_ (.A1(_07819_),
    .A2(_07907_),
    .Z(_07908_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _16029_ (.I(\tt_um_rejunity_sn76489.chan[3].attenuation.control[3] ),
    .ZN(_07909_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _16030_ (.A1(_07909_),
    .A2(_07818_),
    .ZN(_07910_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16031_ (.A1(_07813_),
    .A2(_07822_),
    .ZN(_07911_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16032_ (.A1(_07910_),
    .A2(_07911_),
    .ZN(_07912_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16033_ (.A1(_07820_),
    .A2(_07904_),
    .B(_07912_),
    .ZN(_07913_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _16034_ (.A1(_07908_),
    .A2(_07913_),
    .ZN(_07914_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _16035_ (.A1(_07880_),
    .A2(_07903_),
    .A3(_07914_),
    .Z(_07915_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _16036_ (.I(_07915_),
    .ZN(_07916_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _16037_ (.A1(_07848_),
    .A2(_07863_),
    .Z(_07917_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _16038_ (.A1(_07845_),
    .A2(_07864_),
    .B(_07917_),
    .ZN(_07918_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _16039_ (.A1(_07916_),
    .A2(_07918_),
    .Z(_07919_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _16040_ (.A1(_07873_),
    .A2(_07919_),
    .ZN(_07920_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16041_ (.I(_07868_),
    .Z(_07921_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _16042_ (.A1(\spi_dac_i.spi_dat_buff_1[1] ),
    .A2(_07867_),
    .B1(_07921_),
    .B2(\spi_dac_i.spi_dat_buff_1[2] ),
    .C(_07871_),
    .ZN(_07922_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16043_ (.A1(_07838_),
    .A2(_07920_),
    .B(_07922_),
    .ZN(_00652_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16044_ (.I(_07597_),
    .Z(_07923_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16045_ (.I(_07869_),
    .Z(_07924_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16046_ (.A1(_07873_),
    .A2(_07919_),
    .ZN(_07925_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16047_ (.A1(_07916_),
    .A2(_07918_),
    .B(_07925_),
    .ZN(_07926_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _16048_ (.A1(_07760_),
    .A2(_07875_),
    .ZN(_07927_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16049_ (.A1(_07841_),
    .A2(_07754_),
    .ZN(_07928_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _16050_ (.A1(\tt_um_rejunity_sn76489.chan[2].attenuation.control[2] ),
    .A2(_07927_),
    .B1(_07928_),
    .B2(_07760_),
    .C(_07878_),
    .ZN(_07929_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _16051_ (.I(_07853_),
    .Z(_07930_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _16052_ (.A1(_07784_),
    .A2(_07930_),
    .A3(_07885_),
    .B1(_07887_),
    .B2(_07883_),
    .ZN(_07931_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16053_ (.A1(_07777_),
    .A2(_07890_),
    .ZN(_07932_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _16054_ (.I(_07767_),
    .Z(_07933_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _16055_ (.A1(\tt_um_rejunity_sn76489.chan[1].attenuation.control[2] ),
    .A2(_07933_),
    .A3(_07891_),
    .ZN(_07934_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16056_ (.A1(_07774_),
    .A2(_07778_),
    .B(_07780_),
    .ZN(_07935_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _16057_ (.A1(_07932_),
    .A2(_07934_),
    .A3(_07935_),
    .ZN(_07936_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16058_ (.A1(_07896_),
    .A2(_07902_),
    .B(_07898_),
    .ZN(_07937_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _16059_ (.A1(_07931_),
    .A2(_07936_),
    .A3(_07937_),
    .Z(_07938_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16060_ (.A1(\tt_um_rejunity_sn76489.chan[3].attenuation.control[1] ),
    .A2(_07905_),
    .ZN(_07939_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _16061_ (.I(_07910_),
    .Z(_07940_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _16062_ (.A1(_07823_),
    .A2(_07827_),
    .B(_07817_),
    .C(_07910_),
    .ZN(_07941_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _16063_ (.A1(_07825_),
    .A2(_07823_),
    .B1(_07939_),
    .B2(_07940_),
    .C(_07941_),
    .ZN(_07942_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _16064_ (.A1(_07929_),
    .A2(_07938_),
    .A3(_07942_),
    .ZN(_07943_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _16065_ (.A1(_07903_),
    .A2(_07914_),
    .Z(_07944_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _16066_ (.A1(_07903_),
    .A2(_07914_),
    .Z(_07945_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _16067_ (.A1(_07880_),
    .A2(_07944_),
    .B(_07945_),
    .ZN(_07946_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _16068_ (.A1(_07943_),
    .A2(_07946_),
    .Z(_07947_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _16069_ (.A1(_07926_),
    .A2(_07947_),
    .Z(_07948_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16070_ (.A1(_07926_),
    .A2(_07947_),
    .B(_07721_),
    .ZN(_07949_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16071_ (.A1(\spi_dac_i.spi_dat_buff_1[2] ),
    .A2(_07726_),
    .ZN(_07950_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _16072_ (.A1(_07948_),
    .A2(_07949_),
    .B(_07950_),
    .C(_07869_),
    .ZN(_07951_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16073_ (.A1(\spi_dac_i.spi_dat_buff_1[3] ),
    .A2(_07924_),
    .B(_07951_),
    .ZN(_07952_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16074_ (.A1(_07923_),
    .A2(_07952_),
    .ZN(_00653_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16075_ (.A1(_07943_),
    .A2(_07946_),
    .ZN(_07953_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _16076_ (.A1(_07953_),
    .A2(_07948_),
    .Z(_07954_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16077_ (.I(_07876_),
    .Z(_07955_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16078_ (.A1(_07761_),
    .A2(_07955_),
    .B(_07762_),
    .ZN(_07956_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16079_ (.A1(_07811_),
    .A2(_07906_),
    .ZN(_07957_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _16080_ (.A1(_07811_),
    .A2(_07829_),
    .B(_07957_),
    .ZN(_07958_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _16081_ (.A1(_07930_),
    .A2(_07881_),
    .B(_07804_),
    .ZN(_07959_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _16082_ (.I(_07780_),
    .Z(_07960_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _16083_ (.A1(_07890_),
    .A2(_07778_),
    .ZN(_07961_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16084_ (.A1(_07960_),
    .A2(_07961_),
    .B(_07781_),
    .ZN(_07962_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _16085_ (.A1(_07959_),
    .A2(_07962_),
    .ZN(_07963_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _16086_ (.I(_07931_),
    .ZN(_07964_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16087_ (.A1(_07964_),
    .A2(_07936_),
    .ZN(_07965_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _16088_ (.A1(_07896_),
    .A2(_07902_),
    .A3(_07965_),
    .ZN(_07966_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _16089_ (.A1(_07964_),
    .A2(_07936_),
    .B(_07966_),
    .ZN(_07967_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _16090_ (.A1(_07963_),
    .A2(_07967_),
    .ZN(_07968_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _16091_ (.A1(_07956_),
    .A2(_07958_),
    .A3(_07968_),
    .Z(_07969_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _16092_ (.A1(_07938_),
    .A2(_07942_),
    .Z(_07970_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _16093_ (.A1(_07938_),
    .A2(_07942_),
    .Z(_07971_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _16094_ (.A1(_07929_),
    .A2(_07970_),
    .B(_07971_),
    .ZN(_07972_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _16095_ (.A1(_07954_),
    .A2(_07969_),
    .A3(_07972_),
    .ZN(_07973_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _16096_ (.A1(\spi_dac_i.spi_dat_buff_1[3] ),
    .A2(_07867_),
    .B1(_07921_),
    .B2(\spi_dac_i.spi_dat_buff_1[4] ),
    .C(_07871_),
    .ZN(_07974_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16097_ (.A1(_07838_),
    .A2(_07973_),
    .B(_07974_),
    .ZN(_00654_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16098_ (.A1(_07969_),
    .A2(_07972_),
    .ZN(_07975_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16099_ (.A1(_07969_),
    .A2(_07972_),
    .ZN(_07976_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16100_ (.A1(_07954_),
    .A2(_07975_),
    .B(_07976_),
    .ZN(_07977_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _16101_ (.I(_07956_),
    .ZN(_07978_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16102_ (.A1(_07958_),
    .A2(_07968_),
    .ZN(_07979_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16103_ (.A1(_07958_),
    .A2(_07968_),
    .ZN(_07980_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16104_ (.A1(_07978_),
    .A2(_07979_),
    .B(_07980_),
    .ZN(_07981_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16105_ (.A1(_07749_),
    .A2(_07751_),
    .ZN(_07982_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16106_ (.I(_07747_),
    .Z(_07983_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _16107_ (.A1(_07983_),
    .A2(_07875_),
    .A3(_07955_),
    .ZN(_07984_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _16108_ (.A1(_07982_),
    .A2(_07984_),
    .ZN(_07985_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16109_ (.A1(_07940_),
    .A2(_07907_),
    .ZN(_07986_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _16110_ (.A1(_07824_),
    .A2(_07986_),
    .Z(_07987_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16111_ (.I(_07795_),
    .Z(_07988_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16112_ (.A1(_07988_),
    .A2(_07881_),
    .ZN(_07989_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _16113_ (.A1(_07882_),
    .A2(_07989_),
    .Z(_07990_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _16114_ (.A1(_07800_),
    .A2(_07990_),
    .ZN(_07991_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16115_ (.A1(_07960_),
    .A2(_07892_),
    .ZN(_07992_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _16116_ (.A1(_07776_),
    .A2(_07992_),
    .ZN(_07993_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16117_ (.A1(_07991_),
    .A2(_07993_),
    .ZN(_07994_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _16118_ (.A1(_07991_),
    .A2(_07993_),
    .Z(_07995_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _16119_ (.A1(_07994_),
    .A2(_07995_),
    .Z(_07996_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _16120_ (.A1(_07960_),
    .A2(_07961_),
    .B(_07959_),
    .C(_07781_),
    .ZN(_07997_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16121_ (.A1(_07963_),
    .A2(_07967_),
    .ZN(_07998_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16122_ (.A1(_07997_),
    .A2(_07998_),
    .ZN(_07999_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _16123_ (.A1(_07996_),
    .A2(_07999_),
    .ZN(_08000_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _16124_ (.A1(_07987_),
    .A2(_08000_),
    .Z(_08001_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _16125_ (.A1(_07985_),
    .A2(_08001_),
    .ZN(_08002_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _16126_ (.A1(_07977_),
    .A2(_07981_),
    .A3(_08002_),
    .Z(_08003_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _16127_ (.A1(\spi_dac_i.spi_dat_buff_1[4] ),
    .A2(_07867_),
    .B1(_07921_),
    .B2(\spi_dac_i.spi_dat_buff_1[5] ),
    .C(_03734_),
    .ZN(_08004_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16128_ (.A1(_07743_),
    .A2(_08003_),
    .B(_08004_),
    .ZN(_00655_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _16129_ (.A1(_07981_),
    .A2(_08002_),
    .Z(_08005_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _16130_ (.A1(_07981_),
    .A2(_08002_),
    .Z(_08006_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16131_ (.A1(_07977_),
    .A2(_08005_),
    .B(_08006_),
    .ZN(_08007_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16132_ (.A1(_07757_),
    .A2(_07955_),
    .B(_07843_),
    .ZN(_08008_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16133_ (.A1(_07757_),
    .A2(_07955_),
    .ZN(_08009_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _16134_ (.A1(_07983_),
    .A2(_08008_),
    .B1(_08009_),
    .B2(_07879_),
    .ZN(_08010_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16135_ (.A1(_07825_),
    .A2(_07906_),
    .B(_07846_),
    .ZN(_08011_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16136_ (.A1(_07825_),
    .A2(_07906_),
    .ZN(_08012_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _16137_ (.A1(_07940_),
    .A2(_08011_),
    .B1(_08012_),
    .B2(_07912_),
    .ZN(_08013_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16138_ (.I(_07773_),
    .Z(_08014_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16139_ (.A1(_08014_),
    .A2(_07961_),
    .B(_07858_),
    .ZN(_08015_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16140_ (.A1(_08014_),
    .A2(_07961_),
    .ZN(_08016_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _16141_ (.A1(_07933_),
    .A2(_08015_),
    .B1(_08016_),
    .B2(_07893_),
    .ZN(_08017_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _16142_ (.A1(_07801_),
    .A2(_07786_),
    .B1(_07800_),
    .B2(_07794_),
    .ZN(_08018_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16143_ (.A1(_07792_),
    .A2(_07881_),
    .B(_07886_),
    .ZN(_08019_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16144_ (.A1(_07988_),
    .A2(_08019_),
    .ZN(_08020_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _16145_ (.A1(_07988_),
    .A2(_08018_),
    .B(_08020_),
    .ZN(_08021_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16146_ (.A1(_07996_),
    .A2(_07999_),
    .ZN(_08022_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16147_ (.A1(_07994_),
    .A2(_08022_),
    .ZN(_08023_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _16148_ (.A1(_08017_),
    .A2(_08021_),
    .A3(_08023_),
    .ZN(_08024_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _16149_ (.A1(_08013_),
    .A2(_08024_),
    .ZN(_08025_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _16150_ (.A1(_08010_),
    .A2(_08025_),
    .ZN(_08026_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16151_ (.A1(_07985_),
    .A2(_08001_),
    .ZN(_08027_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16152_ (.A1(_07987_),
    .A2(_08000_),
    .B(_08027_),
    .ZN(_08028_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _16153_ (.A1(_08007_),
    .A2(_08026_),
    .A3(_08028_),
    .ZN(_08029_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _16154_ (.A1(\spi_dac_i.spi_dat_buff_1[5] ),
    .A2(_07729_),
    .B1(_07921_),
    .B2(\spi_dac_i.spi_dat_buff_1[6] ),
    .C(_03734_),
    .ZN(_08030_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16155_ (.A1(_07743_),
    .A2(_08029_),
    .B(_08030_),
    .ZN(_00656_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _16156_ (.A1(_08026_),
    .A2(_08028_),
    .Z(_08031_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _16157_ (.A1(_08026_),
    .A2(_08028_),
    .Z(_08032_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16158_ (.A1(_08007_),
    .A2(_08031_),
    .B(_08032_),
    .ZN(_08033_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _16159_ (.A1(_07983_),
    .A2(_08008_),
    .B1(_08009_),
    .B2(_07879_),
    .C(_08025_),
    .ZN(_08034_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _16160_ (.I(_08034_),
    .ZN(_08035_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _16161_ (.A1(_08013_),
    .A2(_08024_),
    .B(_08035_),
    .ZN(_08036_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _16162_ (.A1(_07759_),
    .A2(_07982_),
    .B1(_07842_),
    .B2(_07877_),
    .ZN(_08037_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16163_ (.A1(\tt_um_rejunity_sn76489.chan[0].attenuation.control[3] ),
    .A2(_07800_),
    .ZN(_08038_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _16164_ (.A1(_07930_),
    .A2(_07850_),
    .A3(_07884_),
    .ZN(_08039_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16165_ (.A1(_08014_),
    .A2(_07892_),
    .B(_07856_),
    .ZN(_08040_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16166_ (.A1(\tt_um_rejunity_sn76489.chan[1].attenuation.control[3] ),
    .A2(_07776_),
    .B(_08040_),
    .ZN(_08041_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16167_ (.A1(_08038_),
    .A2(_08039_),
    .B(_08041_),
    .ZN(_08042_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _16168_ (.A1(_08041_),
    .A2(_08038_),
    .A3(_08039_),
    .Z(_08043_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16169_ (.A1(_08042_),
    .A2(_08043_),
    .ZN(_08044_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _16170_ (.A1(_08017_),
    .A2(_08021_),
    .Z(_08045_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16171_ (.A1(_08017_),
    .A2(_08021_),
    .ZN(_08046_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _16172_ (.I(_08046_),
    .ZN(_08047_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16173_ (.A1(_08045_),
    .A2(_08023_),
    .B(_08047_),
    .ZN(_08048_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _16174_ (.A1(_08044_),
    .A2(_08048_),
    .ZN(_08049_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _16175_ (.A1(_07909_),
    .A2(_07820_),
    .A3(_07823_),
    .B1(_07847_),
    .B2(_07908_),
    .ZN(_08050_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _16176_ (.A1(_08049_),
    .A2(_08050_),
    .Z(_08051_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _16177_ (.A1(_08037_),
    .A2(_08051_),
    .Z(_08052_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _16178_ (.A1(_08033_),
    .A2(_08036_),
    .A3(_08052_),
    .Z(_08053_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _16179_ (.A1(\spi_dac_i.spi_dat_buff_1[6] ),
    .A2(_07729_),
    .B1(_07869_),
    .B2(\spi_dac_i.spi_dat_buff_1[7] ),
    .C(_03734_),
    .ZN(_08054_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16180_ (.A1(_07743_),
    .A2(_08053_),
    .B(_08054_),
    .ZN(_00657_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16181_ (.A1(_08036_),
    .A2(_08052_),
    .ZN(_08055_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16182_ (.A1(_08036_),
    .A2(_08052_),
    .ZN(_08056_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16183_ (.A1(_08033_),
    .A2(_08055_),
    .B(_08056_),
    .ZN(_08057_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _16184_ (.A1(_07761_),
    .A2(_07875_),
    .A3(_07878_),
    .ZN(_08058_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _16185_ (.A1(_07811_),
    .A2(_07904_),
    .A3(_07911_),
    .ZN(_08059_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _16186_ (.I(_07995_),
    .ZN(_08060_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _16187_ (.A1(_07997_),
    .A2(_08060_),
    .B(_08046_),
    .C(_07994_),
    .ZN(_08061_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16188_ (.A1(_08017_),
    .A2(_08021_),
    .ZN(_08062_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16189_ (.A1(_08062_),
    .A2(_08043_),
    .ZN(_08063_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16190_ (.A1(_08061_),
    .A2(_08063_),
    .B(_08042_),
    .ZN(_08064_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _16191_ (.A1(_07933_),
    .A2(_07891_),
    .A3(_07932_),
    .ZN(_08065_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16192_ (.A1(_07882_),
    .A2(_07887_),
    .ZN(_08066_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _16193_ (.A1(_08065_),
    .A2(_08066_),
    .Z(_08067_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _16194_ (.A1(_08064_),
    .A2(_08067_),
    .ZN(_08068_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _16195_ (.A1(_08058_),
    .A2(_08059_),
    .A3(_08068_),
    .ZN(_08069_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _16196_ (.A1(_08049_),
    .A2(_08050_),
    .Z(_08070_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _16197_ (.A1(_08037_),
    .A2(_08051_),
    .B(_08070_),
    .ZN(_08071_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _16198_ (.A1(_08069_),
    .A2(_08071_),
    .Z(_08072_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _16199_ (.A1(_08057_),
    .A2(_08072_),
    .Z(_08073_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16200_ (.A1(_07834_),
    .A2(_08073_),
    .ZN(_08074_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _16201_ (.A1(\spi_dac_i.spi_dat_buff_1[7] ),
    .A2(_07719_),
    .B1(_07870_),
    .B2(\spi_dac_i.spi_dat_buff_1[8] ),
    .C(_07871_),
    .ZN(_08075_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16202_ (.A1(_08074_),
    .A2(_08075_),
    .ZN(_00658_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16203_ (.A1(_08057_),
    .A2(_08072_),
    .ZN(_08076_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _16204_ (.A1(_08069_),
    .A2(_08071_),
    .B(_08076_),
    .ZN(_08077_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16205_ (.A1(_07983_),
    .A2(_07749_),
    .ZN(_08078_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16206_ (.A1(_07940_),
    .A2(_07820_),
    .ZN(_08079_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _16207_ (.A1(_07882_),
    .A2(_07887_),
    .A3(_08065_),
    .ZN(_08080_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16208_ (.A1(_08064_),
    .A2(_08067_),
    .ZN(_08081_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16209_ (.A1(_08080_),
    .A2(_08081_),
    .ZN(_08082_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _16210_ (.A1(_07933_),
    .A2(_07777_),
    .A3(_07930_),
    .A4(_07792_),
    .ZN(_08083_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _16211_ (.A1(_07960_),
    .A2(_08014_),
    .B1(_07988_),
    .B2(_07786_),
    .ZN(_08084_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16212_ (.A1(_08083_),
    .A2(_08084_),
    .ZN(_08085_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _16213_ (.A1(_08082_),
    .A2(_08085_),
    .Z(_08086_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _16214_ (.A1(_08079_),
    .A2(_08086_),
    .ZN(_08087_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _16215_ (.A1(_08078_),
    .A2(_08087_),
    .ZN(_08088_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16216_ (.A1(_08059_),
    .A2(_08068_),
    .ZN(_08089_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16217_ (.A1(_08059_),
    .A2(_08068_),
    .ZN(_08090_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16218_ (.A1(_08058_),
    .A2(_08089_),
    .B(_08090_),
    .ZN(_08091_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _16219_ (.A1(_08088_),
    .A2(_08091_),
    .Z(_08092_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16220_ (.A1(_08077_),
    .A2(_08092_),
    .ZN(_08093_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16221_ (.A1(_08077_),
    .A2(_08092_),
    .ZN(_08094_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16222_ (.A1(_07726_),
    .A2(_08094_),
    .ZN(_08095_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _16223_ (.I(_07727_),
    .Z(_08096_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _16224_ (.A1(\spi_dac_i.spi_dat_buff_1[8] ),
    .A2(_07834_),
    .B1(_08093_),
    .B2(_08095_),
    .C(_08096_),
    .ZN(_08097_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16225_ (.I(_07683_),
    .Z(_08098_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16226_ (.A1(\spi_dac_i.spi_dat_buff_1[9] ),
    .A2(_07924_),
    .B(_08098_),
    .ZN(_08099_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16227_ (.A1(_08097_),
    .A2(_08099_),
    .ZN(_00659_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16228_ (.A1(_08088_),
    .A2(_08091_),
    .ZN(_08100_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16229_ (.A1(_08077_),
    .A2(_08092_),
    .B(_08100_),
    .ZN(_08101_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16230_ (.A1(_08078_),
    .A2(_08087_),
    .ZN(_08102_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16231_ (.A1(_08079_),
    .A2(_08086_),
    .B(_08102_),
    .ZN(_08103_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _16232_ (.A1(_08082_),
    .A2(_08085_),
    .Z(_08104_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16233_ (.A1(_08083_),
    .A2(_08104_),
    .ZN(_08105_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _16234_ (.A1(_08103_),
    .A2(_08105_),
    .Z(_08106_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16235_ (.A1(_08101_),
    .A2(_08106_),
    .B(_07741_),
    .ZN(_08107_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16236_ (.A1(_08101_),
    .A2(_08106_),
    .B(_08107_),
    .ZN(_08108_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _16237_ (.A1(\spi_dac_i.spi_dat_buff_1[9] ),
    .A2(_07834_),
    .B(_08096_),
    .C(_08108_),
    .ZN(_08109_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16238_ (.A1(\spi_dac_i.spi_dat_buff_1[10] ),
    .A2(_07870_),
    .B(_08098_),
    .ZN(_08110_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16239_ (.A1(_08109_),
    .A2(_08110_),
    .ZN(_00660_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16240_ (.A1(_08083_),
    .A2(_08104_),
    .B(_08103_),
    .ZN(_08111_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _16241_ (.A1(\spi_dac_i.spi_dat_buff_1[10] ),
    .A2(_07722_),
    .B1(_08111_),
    .B2(_08107_),
    .ZN(_08112_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16242_ (.A1(\spi_dac_i.spi_dat_buff_1[11] ),
    .A2(_07870_),
    .B(_07700_),
    .ZN(_08113_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16243_ (.A1(_07924_),
    .A2(_08112_),
    .B(_08113_),
    .ZN(_00661_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _16244_ (.A1(\filters.sample_buff[3] ),
    .A2(_07722_),
    .B1(_07728_),
    .B2(\spi_dac_i.spi_dat_buff_0[0] ),
    .ZN(_08114_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16245_ (.A1(_07923_),
    .A2(_08114_),
    .ZN(_00662_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16246_ (.I(_07741_),
    .Z(_08115_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _16247_ (.A1(_07720_),
    .A2(_07717_),
    .ZN(_08116_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16248_ (.I(_08116_),
    .Z(_08117_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _16249_ (.A1(\filters.sample_buff[4] ),
    .A2(_08115_),
    .B1(_08117_),
    .B2(\spi_dac_i.spi_dat_buff_0[0] ),
    .C1(\spi_dac_i.spi_dat_buff_0[1] ),
    .C2(_07728_),
    .ZN(_08118_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16250_ (.A1(_07923_),
    .A2(_08118_),
    .ZN(_00663_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16251_ (.I(_07727_),
    .Z(_08119_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _16252_ (.A1(\filters.sample_buff[5] ),
    .A2(_08115_),
    .B1(_08117_),
    .B2(\spi_dac_i.spi_dat_buff_0[1] ),
    .C1(\spi_dac_i.spi_dat_buff_0[2] ),
    .C2(_08119_),
    .ZN(_08120_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16253_ (.A1(_07923_),
    .A2(_08120_),
    .ZN(_00664_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16254_ (.I(_07597_),
    .Z(_08121_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16255_ (.I(_08116_),
    .Z(_08122_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _16256_ (.A1(\filters.sample_buff[6] ),
    .A2(_08115_),
    .B1(_08122_),
    .B2(\spi_dac_i.spi_dat_buff_0[2] ),
    .C1(\spi_dac_i.spi_dat_buff_0[3] ),
    .C2(_08119_),
    .ZN(_08123_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16257_ (.A1(_08121_),
    .A2(_08123_),
    .ZN(_00665_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _16258_ (.A1(\filters.sample_buff[7] ),
    .A2(_08115_),
    .B1(_08122_),
    .B2(\spi_dac_i.spi_dat_buff_0[3] ),
    .C1(\spi_dac_i.spi_dat_buff_0[4] ),
    .C2(_08119_),
    .ZN(_08124_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16259_ (.A1(_08121_),
    .A2(_08124_),
    .ZN(_00666_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16260_ (.I(_07741_),
    .Z(_08125_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _16261_ (.A1(\filters.sample_buff[8] ),
    .A2(_08125_),
    .B1(_08122_),
    .B2(\spi_dac_i.spi_dat_buff_0[4] ),
    .C1(\spi_dac_i.spi_dat_buff_0[5] ),
    .C2(_08119_),
    .ZN(_08126_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16262_ (.A1(_08121_),
    .A2(_08126_),
    .ZN(_00667_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16263_ (.I(_07727_),
    .Z(_08127_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _16264_ (.A1(\filters.sample_buff[9] ),
    .A2(_08125_),
    .B1(_08122_),
    .B2(\spi_dac_i.spi_dat_buff_0[5] ),
    .C1(\spi_dac_i.spi_dat_buff_0[6] ),
    .C2(_08127_),
    .ZN(_08128_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16265_ (.A1(_08121_),
    .A2(_08128_),
    .ZN(_00668_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _16266_ (.I(_07597_),
    .Z(_08129_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _16267_ (.I(_08116_),
    .Z(_08130_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _16268_ (.A1(\filters.sample_buff[10] ),
    .A2(_08125_),
    .B1(_08130_),
    .B2(\spi_dac_i.spi_dat_buff_0[6] ),
    .C1(\spi_dac_i.spi_dat_buff_0[7] ),
    .C2(_08127_),
    .ZN(_08131_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16269_ (.A1(_08129_),
    .A2(_08131_),
    .ZN(_00669_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _16270_ (.A1(\filters.sample_buff[11] ),
    .A2(_08125_),
    .B1(_08130_),
    .B2(\spi_dac_i.spi_dat_buff_0[7] ),
    .C1(\spi_dac_i.spi_dat_buff_0[8] ),
    .C2(_08127_),
    .ZN(_08132_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16271_ (.A1(_08129_),
    .A2(_08132_),
    .ZN(_00670_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _16272_ (.A1(\filters.sample_buff[12] ),
    .A2(_07742_),
    .B1(_08130_),
    .B2(\spi_dac_i.spi_dat_buff_0[8] ),
    .C1(\spi_dac_i.spi_dat_buff_0[9] ),
    .C2(_08127_),
    .ZN(_08133_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16273_ (.A1(_08129_),
    .A2(_08133_),
    .ZN(_00671_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _16274_ (.A1(\filters.sample_buff[13] ),
    .A2(_07742_),
    .B1(_08130_),
    .B2(\spi_dac_i.spi_dat_buff_0[9] ),
    .C1(\spi_dac_i.spi_dat_buff_0[10] ),
    .C2(_08096_),
    .ZN(_08134_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16275_ (.A1(_08129_),
    .A2(_08134_),
    .ZN(_00672_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _16276_ (.I(_03940_),
    .Z(_08135_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _16277_ (.I(_08135_),
    .Z(_08136_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _16278_ (.A1(\filters.sample_buff[14] ),
    .A2(_07742_),
    .B1(_08116_),
    .B2(\spi_dac_i.spi_dat_buff_0[10] ),
    .C1(\spi_dac_i.spi_dat_buff_0[11] ),
    .C2(_08096_),
    .ZN(_08137_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16279_ (.A1(_08136_),
    .A2(_08137_),
    .ZN(_00673_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16280_ (.A1(net20),
    .A2(_07719_),
    .ZN(_08138_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16281_ (.A1(\spi_dac_i.spi_dat_buff_1[11] ),
    .A2(_08117_),
    .ZN(_08139_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16282_ (.A1(_08138_),
    .A2(_08139_),
    .B(_07740_),
    .ZN(_00674_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16283_ (.A1(net19),
    .A2(_07719_),
    .ZN(_08140_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16284_ (.A1(\spi_dac_i.spi_dat_buff_0[11] ),
    .A2(_08117_),
    .ZN(_08141_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16285_ (.A1(_08140_),
    .A2(_08141_),
    .B(_07740_),
    .ZN(_00675_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16286_ (.A1(_02103_),
    .A2(_07838_),
    .ZN(_00676_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16287_ (.A1(_03738_),
    .A2(_03740_),
    .ZN(_00677_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16288_ (.A1(_02354_),
    .A2(_03741_),
    .ZN(_00678_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _16289_ (.I(\channels.env_counter[3][0] ),
    .Z(_08142_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _16290_ (.I(_08142_),
    .Z(_00679_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _16291_ (.I(\channels.env_counter[3][1] ),
    .Z(_08143_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _16292_ (.I(_08143_),
    .Z(_00680_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _16293_ (.I(\channels.env_counter[3][2] ),
    .Z(_08144_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _16294_ (.I(_08144_),
    .Z(_00681_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _16295_ (.I(\channels.env_counter[3][3] ),
    .Z(_08145_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _16296_ (.I(_08145_),
    .Z(_00682_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _16297_ (.I(\channels.env_counter[3][4] ),
    .Z(_08146_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _16298_ (.I(_08146_),
    .Z(_00683_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _16299_ (.I(\channels.env_counter[3][5] ),
    .Z(_08147_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _16300_ (.I(_08147_),
    .Z(_00684_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _16301_ (.I(\channels.env_counter[3][6] ),
    .Z(_08148_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _16302_ (.I(_08148_),
    .Z(_00685_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _16303_ (.I(\channels.env_counter[3][7] ),
    .Z(_08149_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _16304_ (.I(_08149_),
    .Z(_00686_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _16305_ (.I(\channels.env_counter[3][8] ),
    .Z(_08150_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _16306_ (.I(_08150_),
    .Z(_00687_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _16307_ (.I(\channels.env_counter[3][9] ),
    .Z(_08151_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _16308_ (.I(_08151_),
    .Z(_00688_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _16309_ (.I(\channels.env_counter[3][10] ),
    .Z(_08152_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _16310_ (.I(_08152_),
    .Z(_00689_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _16311_ (.I(\channels.env_counter[3][11] ),
    .Z(_08153_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _16312_ (.I(_08153_),
    .Z(_00690_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _16313_ (.I(\channels.env_counter[3][12] ),
    .Z(_08154_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _16314_ (.I(_08154_),
    .Z(_00691_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _16315_ (.I(\channels.env_counter[3][13] ),
    .Z(_08155_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _16316_ (.I(_08155_),
    .Z(_00692_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _16317_ (.I(\channels.env_counter[3][14] ),
    .Z(_08156_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _16318_ (.I(_08156_),
    .Z(_00693_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16319_ (.A1(_02363_),
    .A2(_03937_),
    .ZN(_08157_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16320_ (.I(_08157_),
    .Z(_08158_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16321_ (.A1(_02363_),
    .A2(_03936_),
    .B(_01821_),
    .ZN(_08159_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16322_ (.I(_08159_),
    .Z(_08160_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16323_ (.A1(\channels.env_vol[1][0] ),
    .A2(_08160_),
    .ZN(_08161_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16324_ (.A1(_03743_),
    .A2(_08158_),
    .B(_08161_),
    .ZN(_00694_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16325_ (.A1(\channels.env_vol[1][1] ),
    .A2(_08160_),
    .ZN(_08162_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16326_ (.A1(_03948_),
    .A2(_08158_),
    .B(_08162_),
    .ZN(_00695_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16327_ (.A1(\channels.env_vol[1][2] ),
    .A2(_08160_),
    .ZN(_08163_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16328_ (.A1(_03954_),
    .A2(_08158_),
    .B(_08163_),
    .ZN(_00696_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16329_ (.A1(\channels.env_vol[1][3] ),
    .A2(_08160_),
    .ZN(_08164_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16330_ (.A1(_03958_),
    .A2(_08158_),
    .B(_08164_),
    .ZN(_00697_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16331_ (.I(_08157_),
    .Z(_08165_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16332_ (.I(_08159_),
    .Z(_08166_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16333_ (.A1(\channels.env_vol[1][4] ),
    .A2(_08166_),
    .ZN(_08167_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16334_ (.A1(_03964_),
    .A2(_08165_),
    .B(_08167_),
    .ZN(_00698_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16335_ (.A1(\channels.env_vol[1][5] ),
    .A2(_08166_),
    .ZN(_08168_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16336_ (.A1(_03974_),
    .A2(_08165_),
    .B(_08168_),
    .ZN(_00699_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16337_ (.A1(\channels.env_vol[1][6] ),
    .A2(_08166_),
    .ZN(_08169_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16338_ (.A1(_03978_),
    .A2(_08165_),
    .B(_08169_),
    .ZN(_00700_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16339_ (.A1(\channels.env_vol[1][7] ),
    .A2(_08166_),
    .ZN(_08170_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16340_ (.A1(_03981_),
    .A2(_08165_),
    .B(_08170_),
    .ZN(_00701_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _16341_ (.A1(_01218_),
    .A2(_01255_),
    .B1(_01258_),
    .B2(\channels.exp_counter[0][0] ),
    .ZN(_08171_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _16342_ (.I(_08171_),
    .ZN(_00702_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _16343_ (.A1(_01225_),
    .A2(_01255_),
    .B1(_01258_),
    .B2(\channels.exp_counter[0][1] ),
    .ZN(_08172_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _16344_ (.I(_08172_),
    .ZN(_00703_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _16345_ (.A1(_01228_),
    .A2(_01317_),
    .B1(_01258_),
    .B2(\channels.exp_counter[0][2] ),
    .ZN(_08173_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _16346_ (.I(_08173_),
    .ZN(_00704_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _16347_ (.A1(_01235_),
    .A2(_01317_),
    .B1(_01334_),
    .B2(\channels.exp_counter[0][3] ),
    .ZN(_08174_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _16348_ (.I(_08174_),
    .ZN(_00705_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _16349_ (.A1(_01238_),
    .A2(_01317_),
    .B1(_01334_),
    .B2(\channels.exp_counter[0][4] ),
    .ZN(_08175_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _16350_ (.I(_08175_),
    .ZN(_00706_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16351_ (.A1(_02356_),
    .A2(_03937_),
    .ZN(_08176_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16352_ (.I(_08176_),
    .Z(_08177_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16353_ (.A1(_02356_),
    .A2(_03936_),
    .B(_01821_),
    .ZN(_08178_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16354_ (.I(_08178_),
    .Z(_08179_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16355_ (.A1(\channels.ch3_env[0] ),
    .A2(_08179_),
    .ZN(_08180_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16356_ (.A1(_03743_),
    .A2(_08177_),
    .B(_08180_),
    .ZN(_00707_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16357_ (.A1(\channels.ch3_env[1] ),
    .A2(_08179_),
    .ZN(_08181_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16358_ (.A1(_03948_),
    .A2(_08177_),
    .B(_08181_),
    .ZN(_00708_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16359_ (.A1(\channels.ch3_env[2] ),
    .A2(_08179_),
    .ZN(_08182_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16360_ (.A1(_03954_),
    .A2(_08177_),
    .B(_08182_),
    .ZN(_00709_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16361_ (.A1(\channels.ch3_env[3] ),
    .A2(_08179_),
    .ZN(_08183_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16362_ (.A1(_03958_),
    .A2(_08177_),
    .B(_08183_),
    .ZN(_00710_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16363_ (.I(_08176_),
    .Z(_08184_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16364_ (.I(_08178_),
    .Z(_08185_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16365_ (.A1(\channels.ch3_env[4] ),
    .A2(_08185_),
    .ZN(_08186_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16366_ (.A1(_03964_),
    .A2(_08184_),
    .B(_08186_),
    .ZN(_00711_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16367_ (.A1(\channels.ch3_env[5] ),
    .A2(_08185_),
    .ZN(_08187_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16368_ (.A1(_03974_),
    .A2(_08184_),
    .B(_08187_),
    .ZN(_00712_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16369_ (.A1(\channels.ch3_env[6] ),
    .A2(_08185_),
    .ZN(_08188_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16370_ (.A1(_03978_),
    .A2(_08184_),
    .B(_08188_),
    .ZN(_00713_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16371_ (.A1(\channels.ch3_env[7] ),
    .A2(_08185_),
    .ZN(_08189_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16372_ (.A1(_03981_),
    .A2(_08184_),
    .B(_08189_),
    .ZN(_00714_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _16373_ (.A1(\tt_um_rejunity_sn76489.noise[0].gen.signal_edge.previous_signal_state_0 ),
    .A2(_02349_),
    .Z(_08190_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16374_ (.I(_08190_),
    .Z(_08191_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16375_ (.I(_08191_),
    .Z(_08192_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16376_ (.A1(\tt_um_rejunity_sn76489.noise[0].gen.lfsr[1] ),
    .A2(_08191_),
    .ZN(_08193_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _16377_ (.A1(\tt_um_rejunity_sn76489.noise[0].gen.restart_noise ),
    .A2(_01042_),
    .Z(_08194_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _16378_ (.I(_08194_),
    .Z(_08195_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _16379_ (.A1(_07809_),
    .A2(_08192_),
    .B(_08193_),
    .C(_08195_),
    .ZN(_00715_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16380_ (.A1(\tt_um_rejunity_sn76489.noise[0].gen.lfsr[1] ),
    .A2(_08192_),
    .ZN(_08196_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _16381_ (.A1(\tt_um_rejunity_sn76489.noise[0].gen.signal_edge.previous_signal_state_0 ),
    .A2(_02349_),
    .ZN(_08197_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16382_ (.I(_08197_),
    .Z(_08198_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16383_ (.A1(\tt_um_rejunity_sn76489.noise[0].gen.lfsr[2] ),
    .A2(_08198_),
    .ZN(_08199_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _16384_ (.I(_08195_),
    .Z(_08200_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16385_ (.A1(_08196_),
    .A2(_08199_),
    .B(_08200_),
    .ZN(_00716_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16386_ (.I(_08191_),
    .Z(_08201_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16387_ (.A1(\tt_um_rejunity_sn76489.noise[0].gen.lfsr[2] ),
    .A2(_08201_),
    .ZN(_08202_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16388_ (.A1(\tt_um_rejunity_sn76489.noise[0].gen.lfsr[3] ),
    .A2(_08198_),
    .ZN(_08203_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16389_ (.A1(_08202_),
    .A2(_08203_),
    .B(_08200_),
    .ZN(_00717_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16390_ (.A1(\tt_um_rejunity_sn76489.noise[0].gen.lfsr[3] ),
    .A2(_08201_),
    .ZN(_08204_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16391_ (.A1(\tt_um_rejunity_sn76489.noise[0].gen.lfsr[4] ),
    .A2(_08198_),
    .ZN(_08205_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16392_ (.A1(_08204_),
    .A2(_08205_),
    .B(_08200_),
    .ZN(_00718_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16393_ (.A1(\tt_um_rejunity_sn76489.noise[0].gen.lfsr[4] ),
    .A2(_08201_),
    .ZN(_08206_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16394_ (.A1(\tt_um_rejunity_sn76489.noise[0].gen.lfsr[5] ),
    .A2(_08198_),
    .ZN(_08207_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16395_ (.A1(_08206_),
    .A2(_08207_),
    .B(_08200_),
    .ZN(_00719_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16396_ (.A1(\tt_um_rejunity_sn76489.noise[0].gen.lfsr[5] ),
    .A2(_08201_),
    .ZN(_08208_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16397_ (.I(_08197_),
    .Z(_08209_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16398_ (.A1(\tt_um_rejunity_sn76489.noise[0].gen.lfsr[6] ),
    .A2(_08209_),
    .ZN(_08210_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _16399_ (.I(_08194_),
    .Z(_08211_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16400_ (.A1(_08208_),
    .A2(_08210_),
    .B(_08211_),
    .ZN(_00720_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _16401_ (.I(_08191_),
    .Z(_08212_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16402_ (.A1(\tt_um_rejunity_sn76489.noise[0].gen.lfsr[6] ),
    .A2(_08212_),
    .ZN(_08213_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16403_ (.A1(\tt_um_rejunity_sn76489.noise[0].gen.lfsr[7] ),
    .A2(_08209_),
    .ZN(_08214_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16404_ (.A1(_08213_),
    .A2(_08214_),
    .B(_08211_),
    .ZN(_00721_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16405_ (.A1(\tt_um_rejunity_sn76489.noise[0].gen.lfsr[7] ),
    .A2(_08212_),
    .ZN(_08215_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16406_ (.A1(\tt_um_rejunity_sn76489.noise[0].gen.lfsr[8] ),
    .A2(_08209_),
    .ZN(_08216_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16407_ (.A1(_08215_),
    .A2(_08216_),
    .B(_08211_),
    .ZN(_00722_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16408_ (.A1(\tt_um_rejunity_sn76489.noise[0].gen.lfsr[8] ),
    .A2(_08212_),
    .ZN(_08217_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16409_ (.A1(\tt_um_rejunity_sn76489.noise[0].gen.lfsr[9] ),
    .A2(_08209_),
    .ZN(_08218_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16410_ (.A1(_08217_),
    .A2(_08218_),
    .B(_08211_),
    .ZN(_00723_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16411_ (.A1(\tt_um_rejunity_sn76489.noise[0].gen.lfsr[9] ),
    .A2(_08212_),
    .ZN(_08219_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16412_ (.I(_08197_),
    .Z(_08220_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16413_ (.A1(\tt_um_rejunity_sn76489.noise[0].gen.lfsr[10] ),
    .A2(_08220_),
    .ZN(_08221_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _16414_ (.I(_08194_),
    .Z(_08222_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16415_ (.A1(_08219_),
    .A2(_08221_),
    .B(_08222_),
    .ZN(_00724_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16416_ (.I(_08190_),
    .Z(_08223_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16417_ (.A1(\tt_um_rejunity_sn76489.noise[0].gen.lfsr[10] ),
    .A2(_08223_),
    .ZN(_08224_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16418_ (.A1(\tt_um_rejunity_sn76489.noise[0].gen.lfsr[11] ),
    .A2(_08220_),
    .ZN(_08225_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16419_ (.A1(_08224_),
    .A2(_08225_),
    .B(_08222_),
    .ZN(_00725_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16420_ (.A1(\tt_um_rejunity_sn76489.noise[0].gen.lfsr[11] ),
    .A2(_08223_),
    .ZN(_08226_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16421_ (.A1(\tt_um_rejunity_sn76489.noise[0].gen.lfsr[12] ),
    .A2(_08220_),
    .ZN(_08227_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16422_ (.A1(_08226_),
    .A2(_08227_),
    .B(_08222_),
    .ZN(_00726_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16423_ (.A1(\tt_um_rejunity_sn76489.noise[0].gen.lfsr[12] ),
    .A2(_08223_),
    .ZN(_08228_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16424_ (.A1(\tt_um_rejunity_sn76489.noise[0].gen.lfsr[13] ),
    .A2(_08220_),
    .ZN(_08229_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16425_ (.A1(_08228_),
    .A2(_08229_),
    .B(_08222_),
    .ZN(_00727_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16426_ (.A1(\tt_um_rejunity_sn76489.noise[0].gen.lfsr[13] ),
    .A2(_08223_),
    .ZN(_08230_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16427_ (.A1(\tt_um_rejunity_sn76489.noise[0].gen.lfsr[14] ),
    .A2(_08197_),
    .ZN(_08231_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16428_ (.A1(_08230_),
    .A2(_08231_),
    .B(_08195_),
    .ZN(_00728_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16429_ (.A1(\tt_um_rejunity_sn76489.control_noise[0][2] ),
    .A2(\tt_um_rejunity_sn76489.noise[0].gen.lfsr[1] ),
    .ZN(_08232_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _16430_ (.A1(_07818_),
    .A2(_08232_),
    .Z(_08233_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16431_ (.A1(\tt_um_rejunity_sn76489.noise[0].gen.lfsr[14] ),
    .A2(_08192_),
    .B(_08195_),
    .ZN(_08234_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16432_ (.A1(_08192_),
    .A2(_08233_),
    .B(_08234_),
    .ZN(_00729_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16433_ (.A1(\tt_um_rejunity_sn76489.clk_counter[4] ),
    .A2(\tt_um_rejunity_sn76489.clk_counter[3] ),
    .ZN(_08235_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _16434_ (.A1(\tt_um_rejunity_sn76489.clk_counter[2] ),
    .A2(\tt_um_rejunity_sn76489.clk_counter[1] ),
    .A3(\tt_um_rejunity_sn76489.clk_counter[0] ),
    .ZN(_08236_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16435_ (.A1(_08235_),
    .A2(_08236_),
    .ZN(_08237_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _16436_ (.I(_08237_),
    .Z(_08238_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _16437_ (.A1(\tt_um_rejunity_sn76489.noise[0].gen.counter[0] ),
    .A2(_08238_),
    .Z(_08239_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16438_ (.A1(_08136_),
    .A2(_08239_),
    .ZN(_00730_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _16439_ (.A1(_08235_),
    .A2(_08236_),
    .Z(_08240_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _16440_ (.I(_08240_),
    .Z(_08241_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16441_ (.I(_08241_),
    .Z(_08242_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _16442_ (.I(_08242_),
    .Z(_08243_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _16443_ (.I(_08243_),
    .Z(_08244_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16444_ (.A1(\tt_um_rejunity_sn76489.noise[0].gen.counter[0] ),
    .A2(_08244_),
    .B(\tt_um_rejunity_sn76489.noise[0].gen.counter[1] ),
    .ZN(_08245_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _16445_ (.A1(\tt_um_rejunity_sn76489.noise[0].gen.counter[1] ),
    .A2(\tt_um_rejunity_sn76489.noise[0].gen.counter[0] ),
    .A3(_08240_),
    .Z(_08246_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _16446_ (.A1(_04101_),
    .A2(_08245_),
    .A3(_08246_),
    .ZN(_00731_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _16447_ (.A1(\tt_um_rejunity_sn76489.noise[0].gen.counter[2] ),
    .A2(_08246_),
    .Z(_08247_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16448_ (.A1(\tt_um_rejunity_sn76489.noise[0].gen.counter[2] ),
    .A2(_08246_),
    .B(_08098_),
    .ZN(_08248_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16449_ (.A1(_08247_),
    .A2(_08248_),
    .ZN(_00732_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _16450_ (.A1(\tt_um_rejunity_sn76489.noise[0].gen.counter[3] ),
    .A2(_08247_),
    .Z(_08249_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16451_ (.A1(\tt_um_rejunity_sn76489.noise[0].gen.counter[3] ),
    .A2(_08247_),
    .B(_08098_),
    .ZN(_08250_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16452_ (.A1(_08249_),
    .A2(_08250_),
    .ZN(_00733_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _16453_ (.A1(\tt_um_rejunity_sn76489.noise[0].gen.counter[4] ),
    .A2(_08249_),
    .Z(_08251_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _16454_ (.I(_07683_),
    .Z(_08252_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16455_ (.A1(\tt_um_rejunity_sn76489.noise[0].gen.counter[4] ),
    .A2(_08249_),
    .B(_08252_),
    .ZN(_08253_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16456_ (.A1(_08251_),
    .A2(_08253_),
    .ZN(_00734_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16457_ (.A1(\tt_um_rejunity_sn76489.noise[0].gen.counter[5] ),
    .A2(_08251_),
    .B(_07700_),
    .ZN(_08254_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16458_ (.A1(\tt_um_rejunity_sn76489.noise[0].gen.counter[5] ),
    .A2(_08251_),
    .B(_08254_),
    .ZN(_00735_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16459_ (.A1(\tt_um_rejunity_sn76489.noise[0].gen.counter[5] ),
    .A2(_08251_),
    .ZN(_08255_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _16460_ (.A1(\tt_um_rejunity_sn76489.noise[0].gen.counter[6] ),
    .A2(_08255_),
    .Z(_08256_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16461_ (.A1(_08136_),
    .A2(_08256_),
    .ZN(_00736_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16462_ (.A1(_08136_),
    .A2(_07924_),
    .ZN(_00737_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16463_ (.I(_08241_),
    .Z(_08257_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _16464_ (.A1(\tt_um_rejunity_sn76489.tone[2].gen.counter[3] ),
    .A2(\tt_um_rejunity_sn76489.tone[2].gen.counter[2] ),
    .A3(\tt_um_rejunity_sn76489.tone[2].gen.counter[1] ),
    .A4(\tt_um_rejunity_sn76489.tone[2].gen.counter[0] ),
    .Z(_08258_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _16465_ (.A1(\tt_um_rejunity_sn76489.tone[2].gen.counter[7] ),
    .A2(\tt_um_rejunity_sn76489.tone[2].gen.counter[6] ),
    .A3(\tt_um_rejunity_sn76489.tone[2].gen.counter[5] ),
    .A4(\tt_um_rejunity_sn76489.tone[2].gen.counter[4] ),
    .Z(_08259_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _16466_ (.A1(\tt_um_rejunity_sn76489.tone[2].gen.counter[9] ),
    .A2(\tt_um_rejunity_sn76489.tone[2].gen.counter[8] ),
    .A3(_08258_),
    .A4(_08259_),
    .ZN(_08260_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _16467_ (.A1(\tt_um_rejunity_sn76489.control_tone_freq[2][0] ),
    .A2(_08260_),
    .B(\tt_um_rejunity_sn76489.tone[2].gen.counter[0] ),
    .ZN(_08261_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16468_ (.A1(_08257_),
    .A2(_08261_),
    .ZN(_08262_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16469_ (.I(_08237_),
    .Z(_08263_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16470_ (.A1(\tt_um_rejunity_sn76489.tone[2].gen.counter[0] ),
    .A2(_08263_),
    .ZN(_08264_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16471_ (.A1(_08262_),
    .A2(_08264_),
    .B(_07740_),
    .ZN(_00738_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16472_ (.I(_08135_),
    .Z(_08265_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _16473_ (.I(\tt_um_rejunity_sn76489.tone[2].gen.counter[1] ),
    .ZN(_08266_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16474_ (.I(_08241_),
    .Z(_08267_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16475_ (.I(_08260_),
    .Z(_08268_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16476_ (.I(_08268_),
    .Z(_08269_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16477_ (.I(_08269_),
    .Z(_08270_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _16478_ (.A1(\tt_um_rejunity_sn76489.control_tone_freq[2][1] ),
    .A2(_08267_),
    .A3(_08270_),
    .ZN(_08271_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16479_ (.A1(_08266_),
    .A2(_08271_),
    .ZN(_08272_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _16480_ (.A1(_08262_),
    .A2(_08272_),
    .Z(_08273_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16481_ (.A1(_08265_),
    .A2(_08273_),
    .ZN(_00739_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16482_ (.I(_08237_),
    .Z(_08274_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16483_ (.A1(\tt_um_rejunity_sn76489.control_tone_freq[2][2] ),
    .A2(_08268_),
    .B(\tt_um_rejunity_sn76489.tone[2].gen.counter[2] ),
    .ZN(_08275_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16484_ (.A1(\tt_um_rejunity_sn76489.control_tone_freq[2][1] ),
    .A2(_08268_),
    .B(\tt_um_rejunity_sn76489.tone[2].gen.counter[1] ),
    .ZN(_08276_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _16485_ (.A1(_08261_),
    .A2(_08275_),
    .A3(_08276_),
    .Z(_08277_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16486_ (.A1(_08261_),
    .A2(_08276_),
    .B(_08275_),
    .ZN(_08278_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _16487_ (.A1(_08274_),
    .A2(_08277_),
    .A3(_08278_),
    .ZN(_08279_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _16488_ (.I(_08241_),
    .Z(_08280_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16489_ (.I(_08280_),
    .Z(_08281_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _16490_ (.I(_08281_),
    .Z(_08282_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16491_ (.A1(\tt_um_rejunity_sn76489.tone[2].gen.counter[2] ),
    .A2(_08282_),
    .B(_08252_),
    .ZN(_08283_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16492_ (.A1(_08279_),
    .A2(_08283_),
    .ZN(_00740_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16493_ (.A1(\tt_um_rejunity_sn76489.control_tone_freq[2][3] ),
    .A2(_08268_),
    .B(\tt_um_rejunity_sn76489.tone[2].gen.counter[3] ),
    .ZN(_08284_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _16494_ (.A1(_08277_),
    .A2(_08284_),
    .Z(_08285_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16495_ (.A1(_08277_),
    .A2(_08284_),
    .B(_08244_),
    .ZN(_08286_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16496_ (.A1(_08285_),
    .A2(_08286_),
    .ZN(_08287_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16497_ (.A1(\tt_um_rejunity_sn76489.tone[2].gen.counter[3] ),
    .A2(_08282_),
    .B(_08252_),
    .ZN(_08288_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16498_ (.A1(_08287_),
    .A2(_08288_),
    .ZN(_00741_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16499_ (.I(_08243_),
    .Z(_08289_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16500_ (.A1(\tt_um_rejunity_sn76489.control_tone_freq[2][4] ),
    .A2(_08269_),
    .B(\tt_um_rejunity_sn76489.tone[2].gen.counter[4] ),
    .ZN(_08290_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _16501_ (.A1(_08285_),
    .A2(_08290_),
    .Z(_08291_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _16502_ (.I(_08257_),
    .Z(_08292_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16503_ (.A1(_08285_),
    .A2(_08290_),
    .B(_08292_),
    .ZN(_08293_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _16504_ (.A1(\tt_um_rejunity_sn76489.tone[2].gen.counter[4] ),
    .A2(_08289_),
    .B1(_08291_),
    .B2(_08293_),
    .ZN(_08294_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16505_ (.A1(_08265_),
    .A2(_08294_),
    .ZN(_00742_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16506_ (.A1(\tt_um_rejunity_sn76489.control_tone_freq[2][5] ),
    .A2(_08269_),
    .B(\tt_um_rejunity_sn76489.tone[2].gen.counter[5] ),
    .ZN(_08295_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _16507_ (.A1(_08291_),
    .A2(_08295_),
    .Z(_08296_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16508_ (.A1(_08291_),
    .A2(_08295_),
    .B(_08292_),
    .ZN(_08297_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _16509_ (.A1(\tt_um_rejunity_sn76489.tone[2].gen.counter[5] ),
    .A2(_08289_),
    .B1(_08296_),
    .B2(_08297_),
    .ZN(_08298_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16510_ (.A1(_08265_),
    .A2(_08298_),
    .ZN(_00743_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16511_ (.A1(\tt_um_rejunity_sn76489.control_tone_freq[2][6] ),
    .A2(_08269_),
    .B(\tt_um_rejunity_sn76489.tone[2].gen.counter[6] ),
    .ZN(_08299_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _16512_ (.A1(_08296_),
    .A2(_08299_),
    .Z(_08300_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _16513_ (.I(_08257_),
    .Z(_08301_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16514_ (.A1(_08296_),
    .A2(_08299_),
    .B(_08301_),
    .ZN(_08302_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _16515_ (.A1(\tt_um_rejunity_sn76489.tone[2].gen.counter[6] ),
    .A2(_08289_),
    .B1(_08300_),
    .B2(_08302_),
    .ZN(_08303_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16516_ (.A1(_08265_),
    .A2(_08303_),
    .ZN(_00744_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16517_ (.A1(\tt_um_rejunity_sn76489.control_tone_freq[2][7] ),
    .A2(_08270_),
    .B(\tt_um_rejunity_sn76489.tone[2].gen.counter[7] ),
    .ZN(_08304_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _16518_ (.A1(_08300_),
    .A2(_08304_),
    .Z(_08305_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16519_ (.A1(_08300_),
    .A2(_08304_),
    .ZN(_08306_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _16520_ (.A1(_08274_),
    .A2(_08305_),
    .A3(_08306_),
    .ZN(_08307_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16521_ (.A1(\tt_um_rejunity_sn76489.tone[2].gen.counter[7] ),
    .A2(_08282_),
    .B(_08252_),
    .ZN(_08308_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16522_ (.A1(_08307_),
    .A2(_08308_),
    .ZN(_00745_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _16523_ (.A1(\tt_um_rejunity_sn76489.control_tone_freq[2][8] ),
    .A2(_08270_),
    .B(\tt_um_rejunity_sn76489.tone[2].gen.counter[8] ),
    .ZN(_08309_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _16524_ (.A1(_08280_),
    .A2(_08305_),
    .A3(_08309_),
    .ZN(_08310_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _16525_ (.A1(_08238_),
    .A2(_08305_),
    .A3(_08309_),
    .ZN(_08311_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16526_ (.A1(\tt_um_rejunity_sn76489.tone[2].gen.counter[8] ),
    .A2(_08263_),
    .B(_08311_),
    .ZN(_08312_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16527_ (.I(_01822_),
    .Z(_08313_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16528_ (.A1(_08310_),
    .A2(_08312_),
    .B(_08313_),
    .ZN(_00746_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16529_ (.I(_08135_),
    .Z(_08314_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _16530_ (.A1(_08242_),
    .A2(_08270_),
    .Z(_08315_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16531_ (.A1(\tt_um_rejunity_sn76489.control_tone_freq[2][9] ),
    .A2(_08315_),
    .B(\tt_um_rejunity_sn76489.tone[2].gen.counter[9] ),
    .ZN(_08316_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _16532_ (.A1(_08310_),
    .A2(_08316_),
    .ZN(_08317_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16533_ (.A1(_08314_),
    .A2(_08317_),
    .ZN(_00747_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _16534_ (.I(_07355_),
    .Z(_08318_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16535_ (.A1(_02347_),
    .A2(_08315_),
    .B(_08318_),
    .ZN(_08319_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16536_ (.A1(_02347_),
    .A2(_08315_),
    .B(_08319_),
    .ZN(_00748_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _16537_ (.A1(\tt_um_rejunity_sn76489.tone[1].gen.counter[3] ),
    .A2(\tt_um_rejunity_sn76489.tone[1].gen.counter[2] ),
    .A3(\tt_um_rejunity_sn76489.tone[1].gen.counter[1] ),
    .A4(\tt_um_rejunity_sn76489.tone[1].gen.counter[0] ),
    .Z(_08320_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _16538_ (.A1(\tt_um_rejunity_sn76489.tone[1].gen.counter[7] ),
    .A2(\tt_um_rejunity_sn76489.tone[1].gen.counter[6] ),
    .A3(\tt_um_rejunity_sn76489.tone[1].gen.counter[5] ),
    .A4(\tt_um_rejunity_sn76489.tone[1].gen.counter[4] ),
    .Z(_08321_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _16539_ (.A1(\tt_um_rejunity_sn76489.tone[1].gen.counter[9] ),
    .A2(\tt_um_rejunity_sn76489.tone[1].gen.counter[8] ),
    .A3(_08320_),
    .A4(_08321_),
    .ZN(_08322_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _16540_ (.A1(\tt_um_rejunity_sn76489.control_tone_freq[1][0] ),
    .A2(_08322_),
    .B(\tt_um_rejunity_sn76489.tone[1].gen.counter[0] ),
    .ZN(_08323_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16541_ (.A1(_08257_),
    .A2(_08323_),
    .ZN(_08324_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16542_ (.A1(\tt_um_rejunity_sn76489.tone[1].gen.counter[0] ),
    .A2(_08263_),
    .ZN(_08325_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16543_ (.A1(_08324_),
    .A2(_08325_),
    .B(_08313_),
    .ZN(_00749_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _16544_ (.I(\tt_um_rejunity_sn76489.tone[1].gen.counter[1] ),
    .ZN(_08326_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16545_ (.I(_08322_),
    .Z(_08327_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16546_ (.I(_08327_),
    .Z(_08328_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16547_ (.I(_08328_),
    .Z(_08329_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _16548_ (.A1(\tt_um_rejunity_sn76489.control_tone_freq[1][1] ),
    .A2(_08267_),
    .A3(_08329_),
    .ZN(_08330_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16549_ (.A1(_08326_),
    .A2(_08330_),
    .ZN(_08331_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _16550_ (.A1(_08324_),
    .A2(_08331_),
    .Z(_08332_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16551_ (.A1(_08314_),
    .A2(_08332_),
    .ZN(_00750_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16552_ (.I(_08237_),
    .Z(_08333_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16553_ (.A1(\tt_um_rejunity_sn76489.control_tone_freq[1][2] ),
    .A2(_08327_),
    .B(\tt_um_rejunity_sn76489.tone[1].gen.counter[2] ),
    .ZN(_08334_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16554_ (.A1(\tt_um_rejunity_sn76489.control_tone_freq[1][1] ),
    .A2(_08327_),
    .B(\tt_um_rejunity_sn76489.tone[1].gen.counter[1] ),
    .ZN(_08335_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _16555_ (.A1(_08323_),
    .A2(_08334_),
    .A3(_08335_),
    .Z(_08336_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16556_ (.A1(_08323_),
    .A2(_08335_),
    .B(_08334_),
    .ZN(_08337_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _16557_ (.A1(_08333_),
    .A2(_08336_),
    .A3(_08337_),
    .ZN(_08338_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16558_ (.I(_01752_),
    .Z(_08339_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16559_ (.A1(\tt_um_rejunity_sn76489.tone[1].gen.counter[2] ),
    .A2(_08282_),
    .B(_08339_),
    .ZN(_08340_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16560_ (.A1(_08338_),
    .A2(_08340_),
    .ZN(_00751_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16561_ (.A1(\tt_um_rejunity_sn76489.control_tone_freq[1][3] ),
    .A2(_08327_),
    .B(\tt_um_rejunity_sn76489.tone[1].gen.counter[3] ),
    .ZN(_08341_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _16562_ (.A1(_08336_),
    .A2(_08341_),
    .Z(_08342_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16563_ (.A1(_08336_),
    .A2(_08341_),
    .B(_08292_),
    .ZN(_08343_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16564_ (.A1(_08342_),
    .A2(_08343_),
    .ZN(_08344_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16565_ (.I(_08243_),
    .Z(_08345_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16566_ (.A1(\tt_um_rejunity_sn76489.tone[1].gen.counter[3] ),
    .A2(_08345_),
    .B(_08339_),
    .ZN(_08346_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16567_ (.A1(_08344_),
    .A2(_08346_),
    .ZN(_00752_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16568_ (.I(_08243_),
    .Z(_08347_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16569_ (.A1(\tt_um_rejunity_sn76489.control_tone_freq[1][4] ),
    .A2(_08328_),
    .B(\tt_um_rejunity_sn76489.tone[1].gen.counter[4] ),
    .ZN(_08348_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _16570_ (.A1(_08342_),
    .A2(_08348_),
    .Z(_08349_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16571_ (.A1(_08342_),
    .A2(_08348_),
    .B(_08301_),
    .ZN(_08350_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _16572_ (.A1(\tt_um_rejunity_sn76489.tone[1].gen.counter[4] ),
    .A2(_08347_),
    .B1(_08349_),
    .B2(_08350_),
    .ZN(_08351_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16573_ (.A1(_08314_),
    .A2(_08351_),
    .ZN(_00753_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16574_ (.A1(\tt_um_rejunity_sn76489.control_tone_freq[1][5] ),
    .A2(_08328_),
    .B(\tt_um_rejunity_sn76489.tone[1].gen.counter[5] ),
    .ZN(_08352_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _16575_ (.A1(_08349_),
    .A2(_08352_),
    .Z(_08353_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16576_ (.A1(_08349_),
    .A2(_08352_),
    .B(_08301_),
    .ZN(_08354_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _16577_ (.A1(\tt_um_rejunity_sn76489.tone[1].gen.counter[5] ),
    .A2(_08347_),
    .B1(_08353_),
    .B2(_08354_),
    .ZN(_08355_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16578_ (.A1(_08314_),
    .A2(_08355_),
    .ZN(_00754_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16579_ (.I(_08135_),
    .Z(_08356_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16580_ (.A1(\tt_um_rejunity_sn76489.control_tone_freq[1][6] ),
    .A2(_08328_),
    .B(\tt_um_rejunity_sn76489.tone[1].gen.counter[6] ),
    .ZN(_08357_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _16581_ (.A1(_08353_),
    .A2(_08357_),
    .Z(_08358_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16582_ (.A1(_08353_),
    .A2(_08357_),
    .B(_08301_),
    .ZN(_08359_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _16583_ (.A1(\tt_um_rejunity_sn76489.tone[1].gen.counter[6] ),
    .A2(_08347_),
    .B1(_08358_),
    .B2(_08359_),
    .ZN(_08360_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16584_ (.A1(_08356_),
    .A2(_08360_),
    .ZN(_00755_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16585_ (.A1(\tt_um_rejunity_sn76489.control_tone_freq[1][7] ),
    .A2(_08329_),
    .B(\tt_um_rejunity_sn76489.tone[1].gen.counter[7] ),
    .ZN(_08361_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _16586_ (.A1(_08358_),
    .A2(_08361_),
    .Z(_08362_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16587_ (.A1(_08358_),
    .A2(_08361_),
    .ZN(_08363_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _16588_ (.A1(_08333_),
    .A2(_08362_),
    .A3(_08363_),
    .ZN(_08364_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16589_ (.A1(\tt_um_rejunity_sn76489.tone[1].gen.counter[7] ),
    .A2(_08345_),
    .B(_08339_),
    .ZN(_08365_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16590_ (.A1(_08364_),
    .A2(_08365_),
    .ZN(_00756_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16591_ (.A1(\tt_um_rejunity_sn76489.control_tone_freq[1][8] ),
    .A2(_08329_),
    .B(\tt_um_rejunity_sn76489.tone[1].gen.counter[8] ),
    .ZN(_08366_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _16592_ (.A1(_08280_),
    .A2(_08362_),
    .A3(_08366_),
    .ZN(_08367_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _16593_ (.A1(_08238_),
    .A2(_08362_),
    .A3(_08366_),
    .ZN(_08368_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16594_ (.A1(\tt_um_rejunity_sn76489.tone[1].gen.counter[8] ),
    .A2(_08274_),
    .B(_08368_),
    .ZN(_08369_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16595_ (.A1(_08367_),
    .A2(_08369_),
    .B(_08313_),
    .ZN(_00757_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _16596_ (.A1(_08242_),
    .A2(_08329_),
    .Z(_08370_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16597_ (.A1(\tt_um_rejunity_sn76489.control_tone_freq[1][9] ),
    .A2(_08370_),
    .B(\tt_um_rejunity_sn76489.tone[1].gen.counter[9] ),
    .ZN(_08371_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _16598_ (.A1(_08367_),
    .A2(_08371_),
    .ZN(_08372_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16599_ (.A1(_08356_),
    .A2(_08372_),
    .ZN(_00758_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16600_ (.A1(\tt_um_rejunity_sn76489.chan[1].attenuation.in ),
    .A2(_08370_),
    .B(_08318_),
    .ZN(_08373_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16601_ (.A1(\tt_um_rejunity_sn76489.chan[1].attenuation.in ),
    .A2(_08370_),
    .B(_08373_),
    .ZN(_00759_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _16602_ (.A1(_01319_),
    .A2(_01587_),
    .Z(_08374_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16603_ (.I(_08374_),
    .Z(_08375_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16604_ (.I(_08375_),
    .Z(_08376_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16605_ (.A1(_01724_),
    .A2(_08374_),
    .ZN(_08377_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16606_ (.I(_08377_),
    .Z(_08378_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16607_ (.I(_08378_),
    .Z(_08379_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _16608_ (.A1(_01580_),
    .A2(_08376_),
    .B1(_08379_),
    .B2(_01595_),
    .ZN(_00760_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _16609_ (.A1(_01598_),
    .A2(_08376_),
    .B1(_08379_),
    .B2(_01601_),
    .ZN(_00761_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _16610_ (.A1(_01608_),
    .A2(_08376_),
    .B1(_08379_),
    .B2(_01612_),
    .ZN(_00762_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _16611_ (.A1(_01615_),
    .A2(_08376_),
    .B1(_08379_),
    .B2(_01617_),
    .ZN(_00763_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16612_ (.I(_08374_),
    .Z(_08380_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16613_ (.I(_08380_),
    .Z(_08381_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16614_ (.I(_08377_),
    .Z(_08382_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16615_ (.I(_08382_),
    .Z(_08383_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _16616_ (.A1(_01620_),
    .A2(_08381_),
    .B1(_08383_),
    .B2(_01622_),
    .ZN(_00764_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _16617_ (.A1(_01625_),
    .A2(_08381_),
    .B1(_08383_),
    .B2(_01629_),
    .ZN(_00765_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _16618_ (.A1(_01632_),
    .A2(_08381_),
    .B1(_08383_),
    .B2(_01635_),
    .ZN(_00766_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _16619_ (.A1(_01638_),
    .A2(_08381_),
    .B1(_08383_),
    .B2(_01640_),
    .ZN(_00767_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16620_ (.I(_08380_),
    .Z(_08384_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16621_ (.I(_08382_),
    .Z(_08385_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _16622_ (.A1(_01645_),
    .A2(_08384_),
    .B1(_08385_),
    .B2(_01647_),
    .ZN(_00768_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _16623_ (.A1(_01650_),
    .A2(_08384_),
    .B1(_08385_),
    .B2(_01653_),
    .ZN(_00769_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _16624_ (.A1(_01657_),
    .A2(_08384_),
    .B1(_08385_),
    .B2(_01660_),
    .ZN(_00770_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _16625_ (.A1(_01663_),
    .A2(_08384_),
    .B1(_08385_),
    .B2(_01665_),
    .ZN(_00771_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16626_ (.I(_08380_),
    .Z(_08386_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16627_ (.I(_08382_),
    .Z(_08387_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _16628_ (.A1(_01668_),
    .A2(_08386_),
    .B1(_08387_),
    .B2(_01670_),
    .ZN(_00772_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _16629_ (.A1(_01673_),
    .A2(_08386_),
    .B1(_08387_),
    .B2(_01676_),
    .ZN(_00773_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _16630_ (.A1(_01681_),
    .A2(_08386_),
    .B1(_08387_),
    .B2(_01684_),
    .ZN(_00774_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _16631_ (.A1(_01689_),
    .A2(_08386_),
    .B1(_08387_),
    .B2(_01691_),
    .ZN(_00775_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16632_ (.I(_08380_),
    .Z(_08388_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16633_ (.I(_08382_),
    .Z(_08389_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _16634_ (.A1(_01694_),
    .A2(_08388_),
    .B1(_08389_),
    .B2(_01695_),
    .ZN(_00776_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _16635_ (.A1(_01698_),
    .A2(_08388_),
    .B1(_08389_),
    .B2(_01573_),
    .ZN(_00777_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _16636_ (.A1(_01577_),
    .A2(_08388_),
    .B1(_08389_),
    .B2(_01702_),
    .ZN(_00778_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _16637_ (.A1(_01705_),
    .A2(_08388_),
    .B1(_08389_),
    .B2(_01707_),
    .ZN(_00779_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _16638_ (.A1(_01710_),
    .A2(_08375_),
    .B1(_08378_),
    .B2(_01712_),
    .ZN(_00780_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _16639_ (.A1(_01715_),
    .A2(_08375_),
    .B1(_08378_),
    .B2(_01717_),
    .ZN(_00781_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _16640_ (.I(\channels.lfsr[0][22] ),
    .ZN(_08390_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _16641_ (.A1(_01720_),
    .A2(_08375_),
    .B1(_08378_),
    .B2(_08390_),
    .ZN(_00782_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _16642_ (.A1(\tt_um_rejunity_sn76489.tone[0].gen.counter[3] ),
    .A2(\tt_um_rejunity_sn76489.tone[0].gen.counter[2] ),
    .A3(\tt_um_rejunity_sn76489.tone[0].gen.counter[1] ),
    .A4(\tt_um_rejunity_sn76489.tone[0].gen.counter[0] ),
    .Z(_08391_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _16643_ (.A1(\tt_um_rejunity_sn76489.tone[0].gen.counter[7] ),
    .A2(\tt_um_rejunity_sn76489.tone[0].gen.counter[6] ),
    .A3(\tt_um_rejunity_sn76489.tone[0].gen.counter[5] ),
    .A4(\tt_um_rejunity_sn76489.tone[0].gen.counter[4] ),
    .Z(_08392_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _16644_ (.A1(\tt_um_rejunity_sn76489.tone[0].gen.counter[9] ),
    .A2(\tt_um_rejunity_sn76489.tone[0].gen.counter[8] ),
    .A3(_08391_),
    .A4(_08392_),
    .ZN(_08393_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _16645_ (.A1(\tt_um_rejunity_sn76489.control_tone_freq[0][0] ),
    .A2(_08393_),
    .B(\tt_um_rejunity_sn76489.tone[0].gen.counter[0] ),
    .ZN(_08394_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16646_ (.A1(_08267_),
    .A2(_08394_),
    .ZN(_08395_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16647_ (.A1(\tt_um_rejunity_sn76489.tone[0].gen.counter[0] ),
    .A2(_08263_),
    .ZN(_08396_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16648_ (.A1(_08395_),
    .A2(_08396_),
    .B(_08313_),
    .ZN(_00783_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _16649_ (.I(\tt_um_rejunity_sn76489.tone[0].gen.counter[1] ),
    .ZN(_08397_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16650_ (.I(_08393_),
    .Z(_08398_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16651_ (.I(_08398_),
    .Z(_08399_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16652_ (.I(_08399_),
    .Z(_08400_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _16653_ (.A1(\tt_um_rejunity_sn76489.control_tone_freq[0][1] ),
    .A2(_08267_),
    .A3(_08400_),
    .ZN(_08401_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16654_ (.A1(_08397_),
    .A2(_08401_),
    .ZN(_08402_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _16655_ (.A1(_08395_),
    .A2(_08402_),
    .Z(_08403_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16656_ (.A1(_08356_),
    .A2(_08403_),
    .ZN(_00784_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16657_ (.A1(\tt_um_rejunity_sn76489.control_tone_freq[0][2] ),
    .A2(_08398_),
    .B(\tt_um_rejunity_sn76489.tone[0].gen.counter[2] ),
    .ZN(_08404_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16658_ (.A1(\tt_um_rejunity_sn76489.control_tone_freq[0][1] ),
    .A2(_08398_),
    .B(\tt_um_rejunity_sn76489.tone[0].gen.counter[1] ),
    .ZN(_08405_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _16659_ (.A1(_08394_),
    .A2(_08404_),
    .A3(_08405_),
    .Z(_08406_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16660_ (.A1(_08394_),
    .A2(_08405_),
    .B(_08404_),
    .ZN(_08407_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _16661_ (.A1(_08333_),
    .A2(_08406_),
    .A3(_08407_),
    .ZN(_08408_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16662_ (.A1(\tt_um_rejunity_sn76489.tone[0].gen.counter[2] ),
    .A2(_08345_),
    .B(_08339_),
    .ZN(_08409_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16663_ (.A1(_08408_),
    .A2(_08409_),
    .ZN(_00785_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16664_ (.A1(\tt_um_rejunity_sn76489.control_tone_freq[0][3] ),
    .A2(_08398_),
    .B(\tt_um_rejunity_sn76489.tone[0].gen.counter[3] ),
    .ZN(_08410_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _16665_ (.A1(_08406_),
    .A2(_08410_),
    .Z(_08411_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16666_ (.A1(_08406_),
    .A2(_08410_),
    .B(_08292_),
    .ZN(_08412_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16667_ (.A1(_08411_),
    .A2(_08412_),
    .ZN(_08413_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16668_ (.A1(\tt_um_rejunity_sn76489.tone[0].gen.counter[3] ),
    .A2(_08345_),
    .B(_01753_),
    .ZN(_08414_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16669_ (.A1(_08413_),
    .A2(_08414_),
    .ZN(_00786_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16670_ (.A1(\tt_um_rejunity_sn76489.control_tone_freq[0][4] ),
    .A2(_08399_),
    .B(\tt_um_rejunity_sn76489.tone[0].gen.counter[4] ),
    .ZN(_08415_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _16671_ (.A1(_08411_),
    .A2(_08415_),
    .Z(_08416_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16672_ (.A1(_08411_),
    .A2(_08415_),
    .B(_08281_),
    .ZN(_08417_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _16673_ (.A1(\tt_um_rejunity_sn76489.tone[0].gen.counter[4] ),
    .A2(_08347_),
    .B1(_08416_),
    .B2(_08417_),
    .ZN(_08418_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16674_ (.A1(_08356_),
    .A2(_08418_),
    .ZN(_00787_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16675_ (.I(_06978_),
    .Z(_08419_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16676_ (.A1(\tt_um_rejunity_sn76489.control_tone_freq[0][5] ),
    .A2(_08399_),
    .B(\tt_um_rejunity_sn76489.tone[0].gen.counter[5] ),
    .ZN(_08420_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _16677_ (.A1(_08416_),
    .A2(_08420_),
    .Z(_08421_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16678_ (.A1(_08416_),
    .A2(_08420_),
    .B(_08281_),
    .ZN(_08422_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _16679_ (.A1(\tt_um_rejunity_sn76489.tone[0].gen.counter[5] ),
    .A2(_08244_),
    .B1(_08421_),
    .B2(_08422_),
    .ZN(_08423_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16680_ (.A1(_08419_),
    .A2(_08423_),
    .ZN(_00788_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16681_ (.A1(\tt_um_rejunity_sn76489.control_tone_freq[0][6] ),
    .A2(_08399_),
    .B(\tt_um_rejunity_sn76489.tone[0].gen.counter[6] ),
    .ZN(_08424_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _16682_ (.A1(_08421_),
    .A2(_08424_),
    .Z(_08425_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16683_ (.A1(_08421_),
    .A2(_08424_),
    .B(_08281_),
    .ZN(_08426_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _16684_ (.A1(\tt_um_rejunity_sn76489.tone[0].gen.counter[6] ),
    .A2(_08244_),
    .B1(_08425_),
    .B2(_08426_),
    .ZN(_08427_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16685_ (.A1(_08419_),
    .A2(_08427_),
    .ZN(_00789_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16686_ (.A1(\tt_um_rejunity_sn76489.control_tone_freq[0][7] ),
    .A2(_08400_),
    .B(\tt_um_rejunity_sn76489.tone[0].gen.counter[7] ),
    .ZN(_08428_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _16687_ (.A1(_08425_),
    .A2(_08428_),
    .Z(_08429_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16688_ (.A1(_08425_),
    .A2(_08428_),
    .ZN(_08430_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _16689_ (.A1(_08333_),
    .A2(_08429_),
    .A3(_08430_),
    .ZN(_08431_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16690_ (.A1(\tt_um_rejunity_sn76489.tone[0].gen.counter[7] ),
    .A2(_08289_),
    .B(_01753_),
    .ZN(_08432_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16691_ (.A1(_08431_),
    .A2(_08432_),
    .ZN(_00790_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _16692_ (.A1(\tt_um_rejunity_sn76489.control_tone_freq[0][8] ),
    .A2(_08400_),
    .B(\tt_um_rejunity_sn76489.tone[0].gen.counter[8] ),
    .ZN(_08433_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _16693_ (.A1(_08280_),
    .A2(_08429_),
    .A3(_08433_),
    .ZN(_08434_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _16694_ (.A1(_08238_),
    .A2(_08429_),
    .A3(_08433_),
    .ZN(_08435_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16695_ (.A1(\tt_um_rejunity_sn76489.tone[0].gen.counter[8] ),
    .A2(_08274_),
    .B(_08435_),
    .ZN(_08436_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16696_ (.A1(_08434_),
    .A2(_08436_),
    .B(_01823_),
    .ZN(_00791_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _16697_ (.A1(_08242_),
    .A2(_08400_),
    .Z(_08437_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16698_ (.A1(\tt_um_rejunity_sn76489.control_tone_freq[0][9] ),
    .A2(_08437_),
    .B(\tt_um_rejunity_sn76489.tone[0].gen.counter[9] ),
    .ZN(_08438_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _16699_ (.A1(_08434_),
    .A2(_08438_),
    .ZN(_08439_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16700_ (.A1(_08419_),
    .A2(_08439_),
    .ZN(_00792_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16701_ (.A1(_07798_),
    .A2(_08437_),
    .B(_08318_),
    .ZN(_08440_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16702_ (.A1(_07798_),
    .A2(_08437_),
    .B(_08440_),
    .ZN(_00793_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _16703_ (.I(\tt_um_rejunity_sn76489.latch_control_reg[2] ),
    .ZN(_08441_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _16704_ (.I(\tt_um_rejunity_sn76489.latch_control_reg[1] ),
    .Z(_08442_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _16705_ (.I(\tt_um_rejunity_sn76489.latch_control_reg[0] ),
    .ZN(_08443_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _16706_ (.A1(_08443_),
    .A2(_01816_),
    .A3(_03494_),
    .ZN(_08444_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _16707_ (.A1(_08441_),
    .A2(_08442_),
    .A3(_08444_),
    .ZN(_08445_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16708_ (.I(_08445_),
    .Z(_08446_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16709_ (.I(_08445_),
    .Z(_08447_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16710_ (.A1(\tt_um_rejunity_sn76489.control_tone_freq[2][4] ),
    .A2(_08447_),
    .B(_08318_),
    .ZN(_08448_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16711_ (.A1(_03710_),
    .A2(_08446_),
    .B(_08448_),
    .ZN(_00794_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _16712_ (.I(_01755_),
    .Z(_08449_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _16713_ (.I(_02100_),
    .Z(_08450_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16714_ (.I(_08450_),
    .Z(_08451_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16715_ (.A1(\tt_um_rejunity_sn76489.control_tone_freq[2][5] ),
    .A2(_08447_),
    .B(_08451_),
    .ZN(_08452_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16716_ (.A1(_08449_),
    .A2(_08446_),
    .B(_08452_),
    .ZN(_00795_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _16717_ (.I(_01765_),
    .Z(_08453_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16718_ (.I(_08445_),
    .Z(_08454_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16719_ (.A1(\tt_um_rejunity_sn76489.control_tone_freq[2][6] ),
    .A2(_08454_),
    .B(_08451_),
    .ZN(_08455_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16720_ (.A1(_08453_),
    .A2(_08446_),
    .B(_08455_),
    .ZN(_00796_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _16721_ (.I(_02298_),
    .Z(_08456_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16722_ (.A1(\tt_um_rejunity_sn76489.control_tone_freq[2][7] ),
    .A2(_08454_),
    .B(_08451_),
    .ZN(_08457_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16723_ (.A1(_08456_),
    .A2(_08446_),
    .B(_08457_),
    .ZN(_00797_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16724_ (.A1(\tt_um_rejunity_sn76489.control_tone_freq[2][8] ),
    .A2(_08454_),
    .B(_08451_),
    .ZN(_08458_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16725_ (.A1(_01800_),
    .A2(_08447_),
    .B(_08458_),
    .ZN(_00798_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16726_ (.I(_08450_),
    .Z(_08459_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16727_ (.A1(\tt_um_rejunity_sn76489.control_tone_freq[2][9] ),
    .A2(_08454_),
    .B(_08459_),
    .ZN(_08460_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16728_ (.A1(_01806_),
    .A2(_08447_),
    .B(_08460_),
    .ZN(_00799_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _16729_ (.I(\tt_um_rejunity_sn76489.latch_control_reg[2] ),
    .Z(_08461_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _16730_ (.I(\tt_um_rejunity_sn76489.latch_control_reg[1] ),
    .ZN(_08462_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _16731_ (.A1(_08461_),
    .A2(_08462_),
    .A3(_08444_),
    .ZN(_08463_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16732_ (.I(_08463_),
    .Z(_08464_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16733_ (.I(_08463_),
    .Z(_08465_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16734_ (.A1(\tt_um_rejunity_sn76489.control_tone_freq[1][4] ),
    .A2(_08465_),
    .B(_08459_),
    .ZN(_08466_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16735_ (.A1(_03710_),
    .A2(_08464_),
    .B(_08466_),
    .ZN(_00800_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16736_ (.A1(\tt_um_rejunity_sn76489.control_tone_freq[1][5] ),
    .A2(_08465_),
    .B(_08459_),
    .ZN(_00860_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16737_ (.A1(_08449_),
    .A2(_08464_),
    .B(_00860_),
    .ZN(_00801_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16738_ (.I(_08463_),
    .Z(_00861_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16739_ (.A1(\tt_um_rejunity_sn76489.control_tone_freq[1][6] ),
    .A2(_00861_),
    .B(_08459_),
    .ZN(_00862_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16740_ (.A1(_08453_),
    .A2(_08464_),
    .B(_00862_),
    .ZN(_00802_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16741_ (.I(_08450_),
    .Z(_00863_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16742_ (.A1(\tt_um_rejunity_sn76489.control_tone_freq[1][7] ),
    .A2(_00861_),
    .B(_00863_),
    .ZN(_00864_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16743_ (.A1(_08456_),
    .A2(_08464_),
    .B(_00864_),
    .ZN(_00803_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16744_ (.A1(\tt_um_rejunity_sn76489.control_tone_freq[1][8] ),
    .A2(_00861_),
    .B(_00863_),
    .ZN(_00865_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16745_ (.A1(_01800_),
    .A2(_08465_),
    .B(_00865_),
    .ZN(_00804_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16746_ (.A1(\tt_um_rejunity_sn76489.control_tone_freq[1][9] ),
    .A2(_00861_),
    .B(_00863_),
    .ZN(_00866_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16747_ (.A1(_01806_),
    .A2(_08465_),
    .B(_00866_),
    .ZN(_00805_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _16748_ (.A1(_08461_),
    .A2(_08442_),
    .A3(_08444_),
    .ZN(_00867_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16749_ (.I(_00867_),
    .Z(_00868_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16750_ (.I(_00867_),
    .Z(_00869_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16751_ (.A1(\tt_um_rejunity_sn76489.control_tone_freq[0][4] ),
    .A2(_00869_),
    .B(_00863_),
    .ZN(_00870_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16752_ (.A1(_03710_),
    .A2(_00868_),
    .B(_00870_),
    .ZN(_00806_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16753_ (.I(_08450_),
    .Z(_00871_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16754_ (.A1(\tt_um_rejunity_sn76489.control_tone_freq[0][5] ),
    .A2(_00869_),
    .B(_00871_),
    .ZN(_00872_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16755_ (.A1(_08449_),
    .A2(_00868_),
    .B(_00872_),
    .ZN(_00807_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16756_ (.I(_00867_),
    .Z(_00873_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16757_ (.A1(\tt_um_rejunity_sn76489.control_tone_freq[0][6] ),
    .A2(_00873_),
    .B(_00871_),
    .ZN(_00874_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16758_ (.A1(_08453_),
    .A2(_00868_),
    .B(_00874_),
    .ZN(_00808_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16759_ (.A1(\tt_um_rejunity_sn76489.control_tone_freq[0][7] ),
    .A2(_00873_),
    .B(_00871_),
    .ZN(_00875_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16760_ (.A1(_08456_),
    .A2(_00868_),
    .B(_00875_),
    .ZN(_00809_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16761_ (.A1(\tt_um_rejunity_sn76489.control_tone_freq[0][8] ),
    .A2(_00873_),
    .B(_00871_),
    .ZN(_00876_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16762_ (.A1(_01800_),
    .A2(_00869_),
    .B(_00876_),
    .ZN(_00810_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _16763_ (.I(_02101_),
    .Z(_00877_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16764_ (.A1(\tt_um_rejunity_sn76489.control_tone_freq[0][9] ),
    .A2(_00873_),
    .B(_00877_),
    .ZN(_00878_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16765_ (.A1(_01806_),
    .A2(_00869_),
    .B(_00878_),
    .ZN(_00811_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16766_ (.I(_03494_),
    .Z(_00879_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16767_ (.A1(\tt_um_rejunity_sn76489.latch_control_reg[0] ),
    .A2(_01816_),
    .ZN(_00880_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16768_ (.A1(_01811_),
    .A2(net15),
    .ZN(_00881_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16769_ (.A1(_03491_),
    .A2(net12),
    .ZN(_00882_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _16770_ (.A1(_08441_),
    .A2(_08462_),
    .A3(_00880_),
    .B1(_00881_),
    .B2(_00882_),
    .ZN(_00883_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _16771_ (.A1(_00879_),
    .A2(_00883_),
    .Z(_00884_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16772_ (.I(_00884_),
    .Z(_00885_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _16773_ (.I(_00884_),
    .Z(_00886_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16774_ (.A1(_03499_),
    .A2(_00886_),
    .ZN(_00887_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _16775_ (.A1(_07826_),
    .A2(_00885_),
    .B(_00887_),
    .C(_02273_),
    .ZN(_00812_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16776_ (.A1(net9),
    .A2(_00886_),
    .ZN(_00888_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16777_ (.I(_02272_),
    .Z(_00889_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _16778_ (.A1(_07821_),
    .A2(_00885_),
    .B(_00888_),
    .C(_00889_),
    .ZN(_00813_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16779_ (.A1(net10),
    .A2(_00886_),
    .ZN(_00890_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _16780_ (.A1(_07817_),
    .A2(_00885_),
    .B(_00890_),
    .C(_00889_),
    .ZN(_00814_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16781_ (.A1(_02098_),
    .A2(_00886_),
    .ZN(_00891_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _16782_ (.A1(_07909_),
    .A2(_00885_),
    .B(_00891_),
    .C(_00889_),
    .ZN(_00815_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _16783_ (.I(\tt_um_rejunity_sn76489.chan[2].attenuation.control[0] ),
    .ZN(_00892_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16784_ (.A1(_01805_),
    .A2(net12),
    .ZN(_00893_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _16785_ (.A1(_08441_),
    .A2(_08442_),
    .A3(_00880_),
    .B1(_00893_),
    .B2(_00881_),
    .ZN(_00894_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _16786_ (.A1(_00879_),
    .A2(_00894_),
    .Z(_00895_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16787_ (.I(_00895_),
    .Z(_00896_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _16788_ (.I(_00895_),
    .Z(_00897_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16789_ (.A1(_03499_),
    .A2(_00897_),
    .ZN(_00898_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _16790_ (.A1(_00892_),
    .A2(_00896_),
    .B(_00898_),
    .C(_00889_),
    .ZN(_00816_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _16791_ (.I(_07841_),
    .ZN(_00899_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16792_ (.A1(net9),
    .A2(_00897_),
    .ZN(_00900_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _16793_ (.I(_02102_),
    .Z(_00901_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _16794_ (.A1(_00899_),
    .A2(_00896_),
    .B(_00900_),
    .C(_00901_),
    .ZN(_00817_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16795_ (.A1(net10),
    .A2(_00897_),
    .ZN(_00902_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _16796_ (.A1(_07755_),
    .A2(_00896_),
    .B(_00902_),
    .C(_00901_),
    .ZN(_00818_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16797_ (.A1(net11),
    .A2(_00897_),
    .ZN(_00903_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _16798_ (.A1(_07759_),
    .A2(_00896_),
    .B(_00903_),
    .C(_00901_),
    .ZN(_00819_));
 gf180mcu_fd_sc_mcu7t5v0__oai33_1 _16799_ (.A1(_03490_),
    .A2(_01817_),
    .A3(_00882_),
    .B1(_00880_),
    .B2(_08462_),
    .B3(_08461_),
    .ZN(_00904_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _16800_ (.A1(_00879_),
    .A2(_00904_),
    .ZN(_00905_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16801_ (.I(_00905_),
    .Z(_00906_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _16802_ (.I(_00905_),
    .Z(_00907_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16803_ (.A1(\tt_um_rejunity_sn76489.chan[1].attenuation.control[0] ),
    .A2(_00907_),
    .ZN(_00908_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _16804_ (.A1(_01741_),
    .A2(_00906_),
    .B(_00908_),
    .C(_00901_),
    .ZN(_00820_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16805_ (.A1(\tt_um_rejunity_sn76489.chan[1].attenuation.control[1] ),
    .A2(_00907_),
    .ZN(_00909_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16806_ (.I(_02102_),
    .Z(_00910_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _16807_ (.A1(_01756_),
    .A2(_00906_),
    .B(_00909_),
    .C(_00910_),
    .ZN(_00821_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16808_ (.A1(\tt_um_rejunity_sn76489.chan[1].attenuation.control[2] ),
    .A2(_00907_),
    .ZN(_00911_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _16809_ (.A1(_08453_),
    .A2(_00906_),
    .B(_00911_),
    .C(_00910_),
    .ZN(_00822_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16810_ (.A1(\tt_um_rejunity_sn76489.chan[1].attenuation.control[3] ),
    .A2(_00907_),
    .ZN(_00912_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _16811_ (.A1(_08456_),
    .A2(_00906_),
    .B(_00912_),
    .C(_00910_),
    .ZN(_00823_));
 gf180mcu_fd_sc_mcu7t5v0__oai33_1 _16812_ (.A1(_08461_),
    .A2(_08442_),
    .A3(_00880_),
    .B1(_00893_),
    .B2(_01817_),
    .B3(_01811_),
    .ZN(_00913_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _16813_ (.A1(_00879_),
    .A2(_00913_),
    .ZN(_00914_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16814_ (.I(_00914_),
    .Z(_00915_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16815_ (.I(_00914_),
    .Z(_00916_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16816_ (.A1(_07801_),
    .A2(_00916_),
    .ZN(_00917_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _16817_ (.A1(_01741_),
    .A2(_00915_),
    .B(_00917_),
    .C(_00910_),
    .ZN(_00824_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16818_ (.A1(\tt_um_rejunity_sn76489.chan[0].attenuation.control[1] ),
    .A2(_00916_),
    .ZN(_00918_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16819_ (.I(_02102_),
    .Z(_00919_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _16820_ (.A1(_01756_),
    .A2(_00915_),
    .B(_00918_),
    .C(_00919_),
    .ZN(_00825_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16821_ (.A1(\tt_um_rejunity_sn76489.chan[0].attenuation.control[2] ),
    .A2(_00916_),
    .ZN(_00920_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _16822_ (.A1(_01766_),
    .A2(_00915_),
    .B(_00920_),
    .C(_00919_),
    .ZN(_00826_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16823_ (.A1(\tt_um_rejunity_sn76489.chan[0].attenuation.control[3] ),
    .A2(_00916_),
    .ZN(_00921_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _16824_ (.A1(_01776_),
    .A2(_00915_),
    .B(_00921_),
    .C(_00919_),
    .ZN(_00827_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _16825_ (.I(_03496_),
    .ZN(_00922_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _16826_ (.A1(_03490_),
    .A2(_00922_),
    .A3(_03519_),
    .ZN(_00923_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16827_ (.A1(\tt_um_rejunity_sn76489.noise[0].gen.restart_noise ),
    .A2(_04158_),
    .ZN(_00924_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16828_ (.A1(_00923_),
    .A2(_00924_),
    .B(_01823_),
    .ZN(_00828_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _16829_ (.I(_03496_),
    .Z(_00925_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16830_ (.A1(_03492_),
    .A2(_00925_),
    .ZN(_00926_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _16831_ (.A1(_08443_),
    .A2(_00925_),
    .B(_00926_),
    .C(_07710_),
    .ZN(_00829_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16832_ (.A1(_03491_),
    .A2(_03496_),
    .ZN(_00927_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _16833_ (.A1(_08462_),
    .A2(_00925_),
    .B(_00927_),
    .C(_04101_),
    .ZN(_00830_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _16834_ (.A1(_08441_),
    .A2(_00925_),
    .B(_03520_),
    .C(_04101_),
    .ZN(_00831_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _16835_ (.I(\tt_um_rejunity_sn76489.clk_counter[0] ),
    .Z(_00928_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16836_ (.A1(_00928_),
    .A2(_03731_),
    .B(_00877_),
    .ZN(_00929_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16837_ (.A1(_00928_),
    .A2(_03732_),
    .B(_00929_),
    .ZN(_00832_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16838_ (.A1(_00928_),
    .A2(_03731_),
    .B(\tt_um_rejunity_sn76489.clk_counter[1] ),
    .ZN(_00930_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _16839_ (.A1(\tt_um_rejunity_sn76489.clk_counter[1] ),
    .A2(_00928_),
    .A3(_03729_),
    .Z(_00931_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _16840_ (.A1(_06917_),
    .A2(_00930_),
    .A3(_00931_),
    .ZN(_00833_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _16841_ (.A1(\tt_um_rejunity_sn76489.clk_counter[2] ),
    .A2(_00931_),
    .Z(_00932_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16842_ (.A1(\tt_um_rejunity_sn76489.clk_counter[2] ),
    .A2(_00931_),
    .B(_01753_),
    .ZN(_00933_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16843_ (.A1(_00932_),
    .A2(_00933_),
    .ZN(_00834_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16844_ (.A1(\tt_um_rejunity_sn76489.clk_counter[3] ),
    .A2(_00932_),
    .B(_00877_),
    .ZN(_00934_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16845_ (.A1(\tt_um_rejunity_sn76489.clk_counter[3] ),
    .A2(_00932_),
    .B(_00934_),
    .ZN(_00835_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16846_ (.A1(\tt_um_rejunity_sn76489.clk_counter[3] ),
    .A2(_00932_),
    .ZN(_00935_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _16847_ (.A1(\tt_um_rejunity_sn76489.clk_counter[4] ),
    .A2(_00935_),
    .Z(_00936_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16848_ (.A1(_08419_),
    .A2(_00936_),
    .ZN(_00836_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _16849_ (.A1(_01581_),
    .A2(_03728_),
    .B(_01087_),
    .ZN(_00937_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16850_ (.I(_00937_),
    .Z(_00938_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16851_ (.I(_00937_),
    .Z(_00939_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _16852_ (.A1(_01583_),
    .A2(_03737_),
    .B(_01092_),
    .C(_01069_),
    .ZN(_00940_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _16853_ (.A1(_02707_),
    .A2(_03742_),
    .ZN(_00941_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _16854_ (.A1(_03096_),
    .A2(_02752_),
    .ZN(_00942_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _16855_ (.A1(_03536_),
    .A2(_03128_),
    .A3(_03131_),
    .A4(_00942_),
    .ZN(_00943_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _16856_ (.A1(_03746_),
    .A2(_00941_),
    .A3(_00943_),
    .Z(_00944_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _16857_ (.A1(_02707_),
    .A2(_03742_),
    .A3(_03128_),
    .A4(_02847_),
    .ZN(_00945_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _16858_ (.A1(_03768_),
    .A2(_03747_),
    .A3(_00942_),
    .A4(_00945_),
    .ZN(_00946_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16859_ (.A1(_00944_),
    .A2(_00946_),
    .ZN(_00947_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16860_ (.A1(_03745_),
    .A2(_03775_),
    .ZN(_00948_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _16861_ (.A1(_03768_),
    .A2(_03971_),
    .A3(_00941_),
    .A4(_00948_),
    .ZN(_00949_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _16862_ (.A1(_03745_),
    .A2(_03752_),
    .A3(_03775_),
    .ZN(_00950_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _16863_ (.A1(_03746_),
    .A2(_00941_),
    .A3(_00950_),
    .ZN(_00951_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _16864_ (.A1(_00947_),
    .A2(_00949_),
    .A3(_00951_),
    .ZN(_00952_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _16865_ (.A1(_01267_),
    .A2(_02455_),
    .B(\channels.clk_div[0] ),
    .C(_01094_),
    .ZN(_00953_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _16866_ (.A1(_03544_),
    .A2(_03755_),
    .A3(_00953_),
    .A4(_00952_),
    .Z(_00954_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _16867_ (.I(_00954_),
    .Z(_00955_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _16868_ (.I(_00955_),
    .ZN(_00956_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _16869_ (.A1(_00940_),
    .A2(_00952_),
    .B1(_00956_),
    .B2(_01183_),
    .ZN(_00957_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16870_ (.A1(_00939_),
    .A2(_00957_),
    .ZN(_00958_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16871_ (.A1(_01180_),
    .A2(_00938_),
    .B(_00958_),
    .ZN(_00837_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16872_ (.A1(_00941_),
    .A2(_00950_),
    .ZN(_00959_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16873_ (.A1(_03746_),
    .A2(_00959_),
    .ZN(_00960_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16874_ (.A1(_00946_),
    .A2(_00960_),
    .B(_00940_),
    .ZN(_00961_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _16875_ (.A1(_01211_),
    .A2(_00955_),
    .B(_00961_),
    .ZN(_00962_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16876_ (.A1(_00939_),
    .A2(_00962_),
    .ZN(_00963_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16877_ (.A1(_01208_),
    .A2(_00938_),
    .B(_00963_),
    .ZN(_00838_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _16878_ (.A1(_00940_),
    .A2(_00954_),
    .ZN(_00964_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16879_ (.A1(_01189_),
    .A2(_00956_),
    .ZN(_00965_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _16880_ (.A1(_00949_),
    .A2(_00964_),
    .B(_00965_),
    .ZN(_00966_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _16881_ (.I0(_00966_),
    .I1(\channels.exp_periods[2][2] ),
    .S(_00937_),
    .Z(_00967_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _16882_ (.I(_00967_),
    .Z(_00839_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16883_ (.A1(_00944_),
    .A2(_00960_),
    .ZN(_00968_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _16884_ (.A1(_01205_),
    .A2(_00955_),
    .B1(_00964_),
    .B2(_00968_),
    .ZN(_00969_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16885_ (.A1(_00939_),
    .A2(_00969_),
    .ZN(_00970_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16886_ (.A1(_01202_),
    .A2(_00938_),
    .B(_00970_),
    .ZN(_00840_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _16887_ (.A1(_01196_),
    .A2(_00955_),
    .B1(_00959_),
    .B2(_00964_),
    .ZN(_00971_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16888_ (.A1(_00939_),
    .A2(_00971_),
    .ZN(_00972_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16889_ (.A1(_01193_),
    .A2(_00938_),
    .B(_00972_),
    .ZN(_00841_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _16890_ (.A1(_01583_),
    .A2(_03739_),
    .ZN(_00973_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _16891_ (.A1(_01724_),
    .A2(_00973_),
    .ZN(_00974_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _16892_ (.I(_00974_),
    .Z(_00975_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _16893_ (.I0(_00957_),
    .I1(\channels.exp_periods[1][0] ),
    .S(_00975_),
    .Z(_00976_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _16894_ (.I(_00976_),
    .Z(_00842_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _16895_ (.I0(_00962_),
    .I1(\channels.exp_periods[1][1] ),
    .S(_00975_),
    .Z(_00977_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _16896_ (.I(_00977_),
    .Z(_00843_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _16897_ (.I0(_00966_),
    .I1(\channels.exp_periods[1][2] ),
    .S(_00975_),
    .Z(_00978_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _16898_ (.I(_00978_),
    .Z(_00844_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _16899_ (.I0(_00969_),
    .I1(\channels.exp_periods[1][3] ),
    .S(_00975_),
    .Z(_00979_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _16900_ (.I(_00979_),
    .Z(_00845_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _16901_ (.I0(_00971_),
    .I1(\channels.exp_periods[1][4] ),
    .S(_00974_),
    .Z(_00980_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _16902_ (.I(_00980_),
    .Z(_00846_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _16903_ (.I(\channels.exp_counter[3][0] ),
    .Z(_00981_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _16904_ (.I(_00981_),
    .Z(_00847_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _16905_ (.I(\channels.exp_counter[3][1] ),
    .Z(_00982_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _16906_ (.I(_00982_),
    .Z(_00848_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _16907_ (.I(\channels.exp_counter[3][2] ),
    .Z(_00983_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _16908_ (.I(_00983_),
    .Z(_00849_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _16909_ (.I(\channels.exp_counter[3][3] ),
    .Z(_00984_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _16910_ (.I(_00984_),
    .Z(_00850_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _16911_ (.I(\channels.exp_counter[3][4] ),
    .Z(_00985_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _16912_ (.I(_00985_),
    .Z(_00851_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _16913_ (.A1(_03744_),
    .A2(_03728_),
    .B(_01043_),
    .ZN(_00986_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _16914_ (.I(_00986_),
    .Z(_00987_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _16915_ (.I0(_00957_),
    .I1(\channels.exp_periods[0][0] ),
    .S(_00987_),
    .Z(_00988_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _16916_ (.I(_00988_),
    .Z(_00852_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _16917_ (.I0(_00962_),
    .I1(\channels.exp_periods[0][1] ),
    .S(_00987_),
    .Z(_00989_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _16918_ (.I(_00989_),
    .Z(_00853_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _16919_ (.I0(_00966_),
    .I1(\channels.exp_periods[0][2] ),
    .S(_00987_),
    .Z(_00990_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _16920_ (.I(_00990_),
    .Z(_00854_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _16921_ (.I0(_00969_),
    .I1(\channels.exp_periods[0][3] ),
    .S(_00987_),
    .Z(_00991_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _16922_ (.I(_00991_),
    .Z(_00855_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _16923_ (.I0(_00971_),
    .I1(\channels.exp_periods[0][4] ),
    .S(_00986_),
    .Z(_00992_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _16924_ (.I(_00992_),
    .Z(_00856_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _16925_ (.A1(_03490_),
    .A2(_00922_),
    .A3(_03519_),
    .Z(_00993_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16926_ (.A1(\tt_um_rejunity_sn76489.control_noise[0][0] ),
    .A2(_00993_),
    .B(_00877_),
    .ZN(_00994_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16927_ (.A1(_01741_),
    .A2(_00993_),
    .B(_00994_),
    .ZN(_00857_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16928_ (.A1(\tt_um_rejunity_sn76489.control_noise[0][1] ),
    .A2(_00993_),
    .B(_02272_),
    .ZN(_00995_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16929_ (.A1(_08449_),
    .A2(_00993_),
    .B(_00995_),
    .ZN(_00858_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16930_ (.A1(\tt_um_rejunity_sn76489.control_noise[0][2] ),
    .A2(_00923_),
    .ZN(_00996_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _16931_ (.A1(_01766_),
    .A2(_00923_),
    .B(_00996_),
    .C(_00919_),
    .ZN(_00859_));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16932_ (.D(_00011_),
    .CLK(clknet_leaf_193_clk),
    .Q(\channels.ring_outs[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16933_ (.D(_00012_),
    .CLK(clknet_leaf_193_clk),
    .Q(\channels.ring_outs[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16934_ (.D(_00013_),
    .CLK(clknet_leaf_215_clk),
    .Q(\channels.lfsr[3][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16935_ (.D(_00014_),
    .CLK(clknet_leaf_216_clk),
    .Q(\channels.lfsr[3][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16936_ (.D(_00015_),
    .CLK(clknet_leaf_216_clk),
    .Q(\channels.lfsr[3][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16937_ (.D(_00016_),
    .CLK(clknet_leaf_217_clk),
    .Q(\channels.lfsr[3][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16938_ (.D(_00017_),
    .CLK(clknet_leaf_220_clk),
    .Q(\channels.lfsr[3][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16939_ (.D(_00018_),
    .CLK(clknet_leaf_220_clk),
    .Q(\channels.lfsr[3][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16940_ (.D(_00019_),
    .CLK(clknet_leaf_220_clk),
    .Q(\channels.lfsr[3][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16941_ (.D(_00020_),
    .CLK(clknet_leaf_221_clk),
    .Q(\channels.lfsr[3][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16942_ (.D(_00021_),
    .CLK(clknet_leaf_221_clk),
    .Q(\channels.lfsr[3][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16943_ (.D(_00022_),
    .CLK(clknet_leaf_226_clk),
    .Q(\channels.lfsr[3][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16944_ (.D(_00023_),
    .CLK(clknet_leaf_227_clk),
    .Q(\channels.lfsr[3][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16945_ (.D(_00024_),
    .CLK(clknet_leaf_227_clk),
    .Q(\channels.lfsr[3][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16946_ (.D(_00025_),
    .CLK(clknet_leaf_236_clk),
    .Q(\channels.lfsr[3][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16947_ (.D(_00026_),
    .CLK(clknet_leaf_238_clk),
    .Q(\channels.lfsr[3][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16948_ (.D(_00027_),
    .CLK(clknet_leaf_239_clk),
    .Q(\channels.lfsr[3][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16949_ (.D(_00028_),
    .CLK(clknet_leaf_238_clk),
    .Q(\channels.lfsr[3][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16950_ (.D(_00029_),
    .CLK(clknet_leaf_239_clk),
    .Q(\channels.lfsr[3][16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16951_ (.D(_00030_),
    .CLK(clknet_leaf_224_clk),
    .Q(\channels.lfsr[3][17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16952_ (.D(_00031_),
    .CLK(clknet_leaf_239_clk),
    .Q(\channels.lfsr[3][18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16953_ (.D(_00032_),
    .CLK(clknet_leaf_239_clk),
    .Q(\channels.lfsr[3][19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16954_ (.D(_00033_),
    .CLK(clknet_leaf_232_clk),
    .Q(\channels.lfsr[3][20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16955_ (.D(_00034_),
    .CLK(clknet_leaf_224_clk),
    .Q(\channels.lfsr[3][21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16956_ (.D(_00035_),
    .CLK(clknet_leaf_212_clk),
    .Q(\channels.lfsr[3][22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16957_ (.D(_00036_),
    .CLK(clknet_leaf_233_clk),
    .Q(\channels.env_vol[3][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16958_ (.D(_00037_),
    .CLK(clknet_5_16__leaf_clk),
    .Q(\channels.env_vol[3][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16959_ (.D(_00038_),
    .CLK(clknet_leaf_232_clk),
    .Q(\channels.env_vol[3][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16960_ (.D(_00039_),
    .CLK(clknet_leaf_211_clk),
    .Q(\channels.env_vol[3][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16961_ (.D(_00040_),
    .CLK(clknet_leaf_213_clk),
    .Q(\channels.env_vol[3][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16962_ (.D(_00041_),
    .CLK(clknet_leaf_233_clk),
    .Q(\channels.env_vol[3][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16963_ (.D(_00042_),
    .CLK(clknet_leaf_211_clk),
    .Q(\channels.env_vol[3][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16964_ (.D(_00043_),
    .CLK(clknet_leaf_211_clk),
    .Q(\channels.env_vol[3][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16965_ (.D(_00044_),
    .CLK(clknet_leaf_194_clk),
    .Q(\channels.exp_counter[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16966_ (.D(_00045_),
    .CLK(clknet_leaf_196_clk),
    .Q(\channels.exp_counter[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16967_ (.D(_00046_),
    .CLK(clknet_leaf_197_clk),
    .Q(\channels.exp_counter[1][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16968_ (.D(_00047_),
    .CLK(clknet_leaf_192_clk),
    .Q(\channels.exp_counter[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16969_ (.D(_00048_),
    .CLK(clknet_leaf_191_clk),
    .Q(\channels.exp_counter[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16970_ (.D(_00049_),
    .CLK(clknet_leaf_193_clk),
    .Q(\channels.exp_counter[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16971_ (.D(_00050_),
    .CLK(clknet_leaf_194_clk),
    .Q(\channels.exp_counter[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16972_ (.D(_00051_),
    .CLK(clknet_5_23__leaf_clk),
    .Q(\channels.exp_counter[2][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16973_ (.D(_00052_),
    .CLK(clknet_leaf_191_clk),
    .Q(\channels.exp_counter[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16974_ (.D(_00053_),
    .CLK(clknet_leaf_191_clk),
    .Q(\channels.exp_counter[2][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16975_ (.D(_00054_),
    .CLK(clknet_leaf_193_clk),
    .Q(\channels.ring_outs[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16976_ (.D(_00055_),
    .CLK(clknet_leaf_187_clk),
    .Q(\channels.accum[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16977_ (.D(_00056_),
    .CLK(clknet_leaf_182_clk),
    .Q(\channels.accum[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16978_ (.D(_00057_),
    .CLK(clknet_leaf_186_clk),
    .Q(\channels.accum[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16979_ (.D(_00058_),
    .CLK(clknet_leaf_180_clk),
    .Q(\channels.accum[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16980_ (.D(_00059_),
    .CLK(clknet_leaf_186_clk),
    .Q(\channels.accum[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16981_ (.D(_00060_),
    .CLK(clknet_leaf_180_clk),
    .Q(\channels.accum[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16982_ (.D(_00061_),
    .CLK(clknet_leaf_188_clk),
    .Q(\channels.accum[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16983_ (.D(_00062_),
    .CLK(clknet_leaf_168_clk),
    .Q(\channels.accum[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16984_ (.D(_00063_),
    .CLK(clknet_leaf_154_clk),
    .Q(\channels.accum[0][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16985_ (.D(_00064_),
    .CLK(clknet_leaf_163_clk),
    .Q(\channels.accum[0][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16986_ (.D(_00065_),
    .CLK(clknet_leaf_152_clk),
    .Q(\channels.accum[0][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16987_ (.D(_00066_),
    .CLK(clknet_leaf_146_clk),
    .Q(\channels.accum[0][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16988_ (.D(_00067_),
    .CLK(clknet_leaf_151_clk),
    .Q(\channels.accum[0][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16989_ (.D(_00068_),
    .CLK(clknet_leaf_164_clk),
    .Q(\channels.accum[0][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16990_ (.D(_00069_),
    .CLK(clknet_leaf_154_clk),
    .Q(\channels.accum[0][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16991_ (.D(_00070_),
    .CLK(clknet_5_28__leaf_clk),
    .Q(\channels.accum[0][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16992_ (.D(_00071_),
    .CLK(clknet_leaf_155_clk),
    .Q(\channels.accum[0][16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16993_ (.D(_00072_),
    .CLK(clknet_leaf_192_clk),
    .Q(\channels.accum[0][17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16994_ (.D(_00073_),
    .CLK(clknet_leaf_156_clk),
    .Q(\channels.accum[0][18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16995_ (.D(_00074_),
    .CLK(clknet_leaf_161_clk),
    .Q(\channels.accum[0][19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16996_ (.D(_00075_),
    .CLK(clknet_leaf_157_clk),
    .Q(\channels.accum[0][20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16997_ (.D(_00076_),
    .CLK(clknet_leaf_189_clk),
    .Q(\channels.accum[0][21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16998_ (.D(_00077_),
    .CLK(clknet_leaf_156_clk),
    .Q(\channels.accum[0][22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16999_ (.D(_00078_),
    .CLK(clknet_leaf_189_clk),
    .Q(\channels.accum[0][23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17000_ (.D(_00079_),
    .CLK(clknet_leaf_212_clk),
    .Q(\channels.lfsr[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17001_ (.D(_00080_),
    .CLK(clknet_leaf_218_clk),
    .Q(\channels.lfsr[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17002_ (.D(_00081_),
    .CLK(clknet_leaf_218_clk),
    .Q(\channels.lfsr[2][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17003_ (.D(_00082_),
    .CLK(clknet_leaf_218_clk),
    .Q(\channels.lfsr[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17004_ (.D(_00083_),
    .CLK(clknet_leaf_219_clk),
    .Q(\channels.lfsr[2][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17005_ (.D(_00084_),
    .CLK(clknet_leaf_219_clk),
    .Q(\channels.lfsr[2][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17006_ (.D(_00085_),
    .CLK(clknet_leaf_224_clk),
    .Q(\channels.lfsr[2][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17007_ (.D(_00086_),
    .CLK(clknet_leaf_222_clk),
    .Q(\channels.lfsr[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17008_ (.D(_00087_),
    .CLK(clknet_leaf_222_clk),
    .Q(\channels.lfsr[2][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17009_ (.D(_00088_),
    .CLK(clknet_leaf_225_clk),
    .Q(\channels.lfsr[2][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17010_ (.D(_00089_),
    .CLK(clknet_leaf_227_clk),
    .Q(\channels.lfsr[2][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17011_ (.D(_00090_),
    .CLK(clknet_leaf_227_clk),
    .Q(\channels.lfsr[2][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17012_ (.D(_00091_),
    .CLK(clknet_leaf_227_clk),
    .Q(\channels.lfsr[2][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17013_ (.D(_00092_),
    .CLK(clknet_leaf_238_clk),
    .Q(\channels.lfsr[2][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17014_ (.D(_00093_),
    .CLK(clknet_leaf_236_clk),
    .Q(\channels.lfsr[2][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17015_ (.D(_00094_),
    .CLK(clknet_leaf_238_clk),
    .Q(\channels.lfsr[2][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17016_ (.D(_00095_),
    .CLK(clknet_5_16__leaf_clk),
    .Q(\channels.lfsr[2][16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17017_ (.D(_00096_),
    .CLK(clknet_leaf_229_clk),
    .Q(\channels.lfsr[2][17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17018_ (.D(_00097_),
    .CLK(clknet_leaf_231_clk),
    .Q(\channels.lfsr[2][18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17019_ (.D(_00098_),
    .CLK(clknet_leaf_235_clk),
    .Q(\channels.lfsr[2][19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17020_ (.D(_00099_),
    .CLK(clknet_leaf_232_clk),
    .Q(\channels.lfsr[2][20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17021_ (.D(_00100_),
    .CLK(clknet_leaf_231_clk),
    .Q(\channels.lfsr[2][21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17022_ (.D(_00101_),
    .CLK(clknet_leaf_212_clk),
    .Q(\channels.lfsr[2][22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17023_ (.D(_00000_),
    .CLK(clknet_leaf_240_clk),
    .Q(\filters.res_lut[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17024_ (.D(_00001_),
    .CLK(clknet_leaf_240_clk),
    .Q(\filters.res_lut[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17025_ (.D(_00002_),
    .CLK(clknet_leaf_240_clk),
    .Q(\filters.res_lut[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17026_ (.D(_00003_),
    .CLK(clknet_leaf_240_clk),
    .Q(\filters.res_lut[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17027_ (.D(_00004_),
    .CLK(clknet_leaf_240_clk),
    .Q(\filters.res_lut[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17028_ (.D(_00005_),
    .CLK(clknet_leaf_240_clk),
    .Q(\filters.res_lut[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17029_ (.D(_00006_),
    .CLK(clknet_leaf_240_clk),
    .Q(\filters.res_lut[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17030_ (.D(_00007_),
    .CLK(clknet_5_18__leaf_clk),
    .Q(\filters.res_lut[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17031_ (.D(_00008_),
    .CLK(clknet_leaf_177_clk),
    .Q(\filters.res_lut[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17032_ (.D(_00102_),
    .CLK(clknet_leaf_213_clk),
    .Q(\channels.lfsr[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17033_ (.D(_00103_),
    .CLK(clknet_leaf_216_clk),
    .Q(\channels.lfsr[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17034_ (.D(_00104_),
    .CLK(clknet_leaf_216_clk),
    .Q(\channels.lfsr[1][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17035_ (.D(_00105_),
    .CLK(clknet_leaf_217_clk),
    .Q(\channels.lfsr[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17036_ (.D(_00106_),
    .CLK(clknet_leaf_221_clk),
    .Q(\channels.lfsr[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17037_ (.D(_00107_),
    .CLK(clknet_leaf_219_clk),
    .Q(\channels.lfsr[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17038_ (.D(_00108_),
    .CLK(clknet_leaf_223_clk),
    .Q(\channels.lfsr[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17039_ (.D(_00109_),
    .CLK(clknet_leaf_223_clk),
    .Q(\channels.lfsr[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17040_ (.D(_00110_),
    .CLK(clknet_leaf_222_clk),
    .Q(\channels.lfsr[1][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17041_ (.D(_00111_),
    .CLK(clknet_leaf_225_clk),
    .Q(\channels.lfsr[1][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17042_ (.D(_00112_),
    .CLK(clknet_leaf_226_clk),
    .Q(\channels.lfsr[1][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17043_ (.D(_00113_),
    .CLK(clknet_leaf_225_clk),
    .Q(\channels.lfsr[1][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17044_ (.D(_00114_),
    .CLK(clknet_leaf_228_clk),
    .Q(\channels.lfsr[1][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17045_ (.D(_00115_),
    .CLK(clknet_leaf_238_clk),
    .Q(\channels.lfsr[1][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17046_ (.D(_00116_),
    .CLK(clknet_leaf_236_clk),
    .Q(\channels.lfsr[1][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17047_ (.D(_00117_),
    .CLK(clknet_leaf_238_clk),
    .Q(\channels.lfsr[1][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17048_ (.D(_00118_),
    .CLK(clknet_5_17__leaf_clk),
    .Q(\channels.lfsr[1][16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17049_ (.D(_00119_),
    .CLK(clknet_leaf_230_clk),
    .Q(\channels.lfsr[1][17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17050_ (.D(_00120_),
    .CLK(clknet_leaf_230_clk),
    .Q(\channels.lfsr[1][18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17051_ (.D(_00121_),
    .CLK(clknet_leaf_230_clk),
    .Q(\channels.lfsr[1][19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17052_ (.D(_00122_),
    .CLK(clknet_leaf_232_clk),
    .Q(\channels.lfsr[1][20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17053_ (.D(_00123_),
    .CLK(clknet_leaf_231_clk),
    .Q(\channels.lfsr[1][21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17054_ (.D(_00124_),
    .CLK(clknet_leaf_212_clk),
    .Q(\channels.lfsr[1][22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17055_ (.D(_00125_),
    .CLK(clknet_leaf_90_clk),
    .Q(\filters.filt_1 ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17056_ (.D(_00126_),
    .CLK(clknet_leaf_89_clk),
    .Q(\filters.filt_2 ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17057_ (.D(_00127_),
    .CLK(clknet_leaf_89_clk),
    .Q(\filters.filt_3 ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17058_ (.D(_00128_),
    .CLK(clknet_leaf_76_clk),
    .Q(\filters.res_filt[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17059_ (.D(_00129_),
    .CLK(clknet_leaf_94_clk),
    .Q(\filters.res_filt[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17060_ (.D(_00130_),
    .CLK(clknet_leaf_178_clk),
    .Q(\filters.res_filt[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17061_ (.D(_00131_),
    .CLK(clknet_leaf_176_clk),
    .Q(\filters.res_filt[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17062_ (.D(_00132_),
    .CLK(clknet_leaf_177_clk),
    .Q(\filters.res_filt[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17063_ (.D(_00133_),
    .CLK(clknet_leaf_105_clk),
    .Q(\filters.mode_vol[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17064_ (.D(_00134_),
    .CLK(clknet_leaf_105_clk),
    .Q(\filters.mode_vol[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17065_ (.D(_00135_),
    .CLK(clknet_leaf_106_clk),
    .Q(\filters.mode_vol[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17066_ (.D(_00136_),
    .CLK(clknet_leaf_106_clk),
    .Q(\filters.mode_vol[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17067_ (.D(_00137_),
    .CLK(clknet_leaf_104_clk),
    .Q(\filters.lp ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17068_ (.D(_00138_),
    .CLK(clknet_leaf_99_clk),
    .Q(\filters.bp ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17069_ (.D(_00139_),
    .CLK(clknet_leaf_98_clk),
    .Q(\filters.hp ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17070_ (.D(_00140_),
    .CLK(clknet_leaf_99_clk),
    .Q(\filters.mode_vol[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17071_ (.D(_00141_),
    .CLK(clknet_leaf_119_clk),
    .Q(net22));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17072_ (.D(_00142_),
    .CLK(clknet_leaf_113_clk),
    .Q(net23));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17073_ (.D(_00143_),
    .CLK(clknet_leaf_119_clk),
    .Q(net24));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17074_ (.D(_00144_),
    .CLK(clknet_leaf_119_clk),
    .Q(net25));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17075_ (.D(_00145_),
    .CLK(clknet_leaf_119_clk),
    .Q(net26));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17076_ (.D(_00146_),
    .CLK(clknet_leaf_119_clk),
    .Q(net27));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17077_ (.D(_00147_),
    .CLK(clknet_leaf_125_clk),
    .Q(net28));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17078_ (.D(_00148_),
    .CLK(clknet_leaf_119_clk),
    .Q(net29));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17079_ (.D(_00149_),
    .CLK(clknet_leaf_107_clk),
    .Q(\channels.freq1[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17080_ (.D(_00150_),
    .CLK(clknet_leaf_107_clk),
    .Q(\channels.freq1[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17081_ (.D(_00151_),
    .CLK(clknet_leaf_107_clk),
    .Q(\channels.freq1[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17082_ (.D(_00152_),
    .CLK(clknet_leaf_106_clk),
    .Q(\channels.freq1[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17083_ (.D(_00153_),
    .CLK(clknet_leaf_109_clk),
    .Q(\channels.freq1[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17084_ (.D(_00154_),
    .CLK(clknet_leaf_108_clk),
    .Q(\channels.freq1[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17085_ (.D(_00155_),
    .CLK(clknet_leaf_109_clk),
    .Q(\channels.freq1[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17086_ (.D(_00156_),
    .CLK(clknet_leaf_109_clk),
    .Q(\channels.freq1[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17087_ (.D(_00157_),
    .CLK(clknet_leaf_107_clk),
    .Q(\channels.pw1[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17088_ (.D(_00158_),
    .CLK(clknet_leaf_112_clk),
    .Q(\channels.pw1[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17089_ (.D(_00159_),
    .CLK(clknet_leaf_107_clk),
    .Q(\channels.pw1[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17090_ (.D(_00160_),
    .CLK(clknet_leaf_113_clk),
    .Q(\channels.pw1[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17091_ (.D(_00161_),
    .CLK(clknet_leaf_110_clk),
    .Q(\channels.ctrl_reg1[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17092_ (.D(_00162_),
    .CLK(clknet_leaf_110_clk),
    .Q(\channels.ctrl_reg1[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17093_ (.D(_00163_),
    .CLK(clknet_leaf_110_clk),
    .Q(\channels.ctrl_reg1[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17094_ (.D(_00164_),
    .CLK(clknet_leaf_110_clk),
    .Q(\channels.ctrl_reg1[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17095_ (.D(_00165_),
    .CLK(clknet_leaf_104_clk),
    .Q(\channels.ctrl_reg1[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17096_ (.D(_00166_),
    .CLK(clknet_leaf_99_clk),
    .Q(\channels.ctrl_reg1[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17097_ (.D(_00167_),
    .CLK(clknet_leaf_99_clk),
    .Q(\channels.ctrl_reg1[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17098_ (.D(_00168_),
    .CLK(clknet_leaf_98_clk),
    .Q(\channels.ctrl_reg1[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17099_ (.D(_00169_),
    .CLK(clknet_leaf_111_clk),
    .Q(\channels.atk_dec1[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17100_ (.D(_00170_),
    .CLK(clknet_leaf_111_clk),
    .Q(\channels.atk_dec1[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17101_ (.D(_00171_),
    .CLK(clknet_leaf_112_clk),
    .Q(\channels.atk_dec1[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17102_ (.D(_00172_),
    .CLK(clknet_leaf_111_clk),
    .Q(\channels.atk_dec1[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17103_ (.D(_00173_),
    .CLK(clknet_leaf_110_clk),
    .Q(\channels.atk_dec1[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17104_ (.D(_00174_),
    .CLK(clknet_leaf_109_clk),
    .Q(\channels.atk_dec1[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17105_ (.D(_00175_),
    .CLK(clknet_leaf_108_clk),
    .Q(\channels.atk_dec1[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17106_ (.D(_00176_),
    .CLK(clknet_leaf_109_clk),
    .Q(\channels.atk_dec1[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17107_ (.D(_00177_),
    .CLK(clknet_leaf_112_clk),
    .Q(\channels.sus_rel1[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17108_ (.D(_00178_),
    .CLK(clknet_leaf_111_clk),
    .Q(\channels.sus_rel1[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17109_ (.D(_00179_),
    .CLK(clknet_leaf_114_clk),
    .Q(\channels.sus_rel1[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17110_ (.D(_00180_),
    .CLK(clknet_leaf_114_clk),
    .Q(\channels.sus_rel1[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17111_ (.D(_00181_),
    .CLK(clknet_leaf_114_clk),
    .Q(\channels.sus_rel1[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17112_ (.D(_00182_),
    .CLK(clknet_leaf_116_clk),
    .Q(\channels.sus_rel1[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17113_ (.D(_00183_),
    .CLK(clknet_leaf_116_clk),
    .Q(\channels.sus_rel1[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17114_ (.D(_00184_),
    .CLK(clknet_leaf_116_clk),
    .Q(\channels.sus_rel1[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17115_ (.D(_00185_),
    .CLK(clknet_leaf_111_clk),
    .Q(\channels.freq2[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17116_ (.D(_00186_),
    .CLK(clknet_leaf_111_clk),
    .Q(\channels.freq2[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17117_ (.D(_00187_),
    .CLK(clknet_leaf_115_clk),
    .Q(\channels.freq2[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17118_ (.D(_00188_),
    .CLK(clknet_leaf_114_clk),
    .Q(\channels.freq2[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17119_ (.D(_00189_),
    .CLK(clknet_leaf_115_clk),
    .Q(\channels.freq2[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17120_ (.D(_00190_),
    .CLK(clknet_leaf_115_clk),
    .Q(\channels.freq2[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17121_ (.D(_00191_),
    .CLK(clknet_leaf_116_clk),
    .Q(\channels.freq2[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17122_ (.D(_00192_),
    .CLK(clknet_leaf_116_clk),
    .Q(\channels.freq2[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17123_ (.D(_00193_),
    .CLK(clknet_leaf_119_clk),
    .Q(\channels.pw2[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17124_ (.D(_00194_),
    .CLK(clknet_leaf_118_clk),
    .Q(\channels.pw2[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17125_ (.D(_00195_),
    .CLK(clknet_leaf_117_clk),
    .Q(\channels.pw2[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17126_ (.D(_00196_),
    .CLK(clknet_leaf_113_clk),
    .Q(\channels.pw2[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17127_ (.D(_00197_),
    .CLK(clknet_leaf_127_clk),
    .Q(\channels.ctrl_reg2[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17128_ (.D(_00198_),
    .CLK(clknet_5_27__leaf_clk),
    .Q(\channels.ctrl_reg2[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17129_ (.D(_00199_),
    .CLK(clknet_leaf_118_clk),
    .Q(\channels.ctrl_reg2[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17130_ (.D(_00200_),
    .CLK(clknet_leaf_117_clk),
    .Q(\channels.ctrl_reg2[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17131_ (.D(_00201_),
    .CLK(clknet_leaf_127_clk),
    .Q(\channels.ctrl_reg2[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17132_ (.D(_00202_),
    .CLK(clknet_leaf_117_clk),
    .Q(\channels.ctrl_reg2[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17133_ (.D(_00203_),
    .CLK(clknet_leaf_117_clk),
    .Q(\channels.ctrl_reg2[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17134_ (.D(_00204_),
    .CLK(clknet_leaf_127_clk),
    .Q(\channels.ctrl_reg2[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17135_ (.D(_00205_),
    .CLK(clknet_leaf_128_clk),
    .Q(\channels.atk_dec2[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17136_ (.D(_00206_),
    .CLK(clknet_leaf_124_clk),
    .Q(\channels.atk_dec2[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17137_ (.D(_00207_),
    .CLK(clknet_leaf_127_clk),
    .Q(\channels.atk_dec2[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17138_ (.D(_00208_),
    .CLK(clknet_leaf_124_clk),
    .Q(\channels.atk_dec2[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17139_ (.D(_00209_),
    .CLK(clknet_leaf_127_clk),
    .Q(\channels.atk_dec2[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17140_ (.D(_00210_),
    .CLK(clknet_leaf_128_clk),
    .Q(\channels.atk_dec2[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17141_ (.D(_00211_),
    .CLK(clknet_leaf_127_clk),
    .Q(\channels.atk_dec2[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17142_ (.D(_00212_),
    .CLK(clknet_leaf_128_clk),
    .Q(\channels.atk_dec2[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17143_ (.D(_00213_),
    .CLK(clknet_leaf_128_clk),
    .Q(\channels.sus_rel2[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17144_ (.D(_00214_),
    .CLK(clknet_leaf_123_clk),
    .Q(\channels.sus_rel2[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17145_ (.D(_00215_),
    .CLK(clknet_leaf_124_clk),
    .Q(\channels.sus_rel2[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17146_ (.D(_00216_),
    .CLK(clknet_leaf_123_clk),
    .Q(\channels.sus_rel2[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17147_ (.D(_00217_),
    .CLK(clknet_leaf_144_clk),
    .Q(\channels.sus_rel2[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17148_ (.D(_00218_),
    .CLK(clknet_leaf_145_clk),
    .Q(\channels.sus_rel2[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17149_ (.D(_00219_),
    .CLK(clknet_leaf_142_clk),
    .Q(\channels.sus_rel2[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17150_ (.D(_00220_),
    .CLK(clknet_leaf_142_clk),
    .Q(\channels.sus_rel2[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17151_ (.D(_00221_),
    .CLK(clknet_leaf_143_clk),
    .Q(\channels.freq3[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17152_ (.D(_00222_),
    .CLK(clknet_leaf_143_clk),
    .Q(\channels.freq3[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17153_ (.D(_00223_),
    .CLK(clknet_leaf_122_clk),
    .Q(\channels.freq3[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17154_ (.D(_00224_),
    .CLK(clknet_leaf_141_clk),
    .Q(\channels.freq3[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17155_ (.D(_00225_),
    .CLK(clknet_leaf_141_clk),
    .Q(\channels.freq3[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17156_ (.D(_00226_),
    .CLK(clknet_leaf_141_clk),
    .Q(\channels.freq3[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17157_ (.D(_00227_),
    .CLK(clknet_leaf_142_clk),
    .Q(\channels.freq3[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17158_ (.D(_00228_),
    .CLK(clknet_leaf_142_clk),
    .Q(\channels.freq3[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17159_ (.D(_00229_),
    .CLK(clknet_leaf_121_clk),
    .Q(\channels.pw3[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17160_ (.D(_00230_),
    .CLK(clknet_leaf_166_clk),
    .Q(\channels.pw3[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17161_ (.D(_00231_),
    .CLK(clknet_leaf_121_clk),
    .Q(\channels.pw3[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17162_ (.D(_00232_),
    .CLK(clknet_5_26__leaf_clk),
    .Q(\channels.pw3[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17163_ (.D(_00233_),
    .CLK(clknet_leaf_144_clk),
    .Q(\channels.ctrl_reg3[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17164_ (.D(_00234_),
    .CLK(clknet_leaf_144_clk),
    .Q(\channels.ctrl_reg3[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17165_ (.D(_00235_),
    .CLK(clknet_leaf_144_clk),
    .Q(\channels.ctrl_reg3[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17166_ (.D(_00236_),
    .CLK(clknet_leaf_143_clk),
    .Q(\channels.ctrl_reg3[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17167_ (.D(_00237_),
    .CLK(clknet_leaf_146_clk),
    .Q(\channels.ctrl_reg3[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17168_ (.D(_00238_),
    .CLK(clknet_leaf_145_clk),
    .Q(\channels.ctrl_reg3[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17169_ (.D(_00239_),
    .CLK(clknet_leaf_145_clk),
    .Q(\channels.ctrl_reg3[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17170_ (.D(_00240_),
    .CLK(clknet_leaf_144_clk),
    .Q(\channels.ctrl_reg3[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17171_ (.D(_00241_),
    .CLK(clknet_leaf_125_clk),
    .Q(\channels.atk_dec3[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17172_ (.D(_00242_),
    .CLK(clknet_leaf_125_clk),
    .Q(\channels.atk_dec3[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17173_ (.D(_00243_),
    .CLK(clknet_leaf_125_clk),
    .Q(\channels.atk_dec3[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17174_ (.D(_00244_),
    .CLK(clknet_leaf_118_clk),
    .Q(\channels.atk_dec3[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17175_ (.D(_00245_),
    .CLK(clknet_leaf_141_clk),
    .Q(\channels.atk_dec3[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17176_ (.D(_00246_),
    .CLK(clknet_leaf_123_clk),
    .Q(\channels.atk_dec3[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17177_ (.D(_00247_),
    .CLK(clknet_leaf_123_clk),
    .Q(\channels.atk_dec3[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17178_ (.D(_00248_),
    .CLK(clknet_leaf_122_clk),
    .Q(\channels.atk_dec3[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17179_ (.D(_00249_),
    .CLK(clknet_leaf_76_clk),
    .Q(\channels.sus_rel3[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17180_ (.D(_00250_),
    .CLK(clknet_leaf_76_clk),
    .Q(\channels.sus_rel3[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17181_ (.D(_00251_),
    .CLK(clknet_leaf_72_clk),
    .Q(\channels.sus_rel3[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17182_ (.D(_00252_),
    .CLK(clknet_leaf_106_clk),
    .Q(\channels.sus_rel3[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17183_ (.D(_00253_),
    .CLK(clknet_leaf_104_clk),
    .Q(\channels.sus_rel3[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17184_ (.D(_00254_),
    .CLK(clknet_leaf_104_clk),
    .Q(\channels.sus_rel3[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17185_ (.D(_00255_),
    .CLK(clknet_leaf_105_clk),
    .Q(\channels.sus_rel3[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17186_ (.D(_00256_),
    .CLK(clknet_leaf_105_clk),
    .Q(\channels.sus_rel3[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17187_ (.D(_00257_),
    .CLK(clknet_leaf_78_clk),
    .Q(\filters.cutoff_lut[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17188_ (.D(_00258_),
    .CLK(clknet_leaf_79_clk),
    .Q(\filters.cutoff_lut[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17189_ (.D(_00259_),
    .CLK(clknet_leaf_78_clk),
    .Q(\filters.cutoff_lut[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17190_ (.D(_00260_),
    .CLK(clknet_leaf_78_clk),
    .Q(\filters.cutoff_lut[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17191_ (.D(_00261_),
    .CLK(clknet_leaf_89_clk),
    .Q(\filters.cutoff_lut[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17192_ (.D(_00262_),
    .CLK(clknet_leaf_89_clk),
    .Q(\filters.cutoff_lut[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17193_ (.D(_00263_),
    .CLK(clknet_leaf_89_clk),
    .Q(\filters.cutoff_lut[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17194_ (.D(_00264_),
    .CLK(clknet_leaf_89_clk),
    .Q(\filters.cutoff_lut[16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17195_ (.D(_00265_),
    .CLK(clknet_leaf_53_clk),
    .Q(\tt_um_rejunity_sn76489.noise[0].gen.signal_edge.previous_signal_state_0 ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17196_ (.D(_00266_),
    .CLK(clknet_leaf_78_clk),
    .Q(\clk_trg[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17197_ (.D(_00267_),
    .CLK(clknet_leaf_79_clk),
    .Q(\clk_trg[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17198_ (.D(_00268_),
    .CLK(clknet_leaf_168_clk),
    .Q(\channels.sync_outs[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17199_ (.D(_00269_),
    .CLK(clknet_leaf_168_clk),
    .Q(\channels.sync_outs[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17200_ (.D(_00270_),
    .CLK(clknet_leaf_168_clk),
    .Q(\channels.sync_outs[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17201_ (.D(_00271_),
    .CLK(clknet_leaf_169_clk),
    .Q(\channels.sample3[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17202_ (.D(_00272_),
    .CLK(clknet_leaf_179_clk),
    .Q(\channels.sample3[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17203_ (.D(_00273_),
    .CLK(clknet_leaf_179_clk),
    .Q(\channels.sample3[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17204_ (.D(_00274_),
    .CLK(clknet_leaf_174_clk),
    .Q(\channels.sample3[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17205_ (.D(_00275_),
    .CLK(clknet_leaf_174_clk),
    .Q(\channels.sample3[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17206_ (.D(_00276_),
    .CLK(clknet_leaf_174_clk),
    .Q(\channels.sample3[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17207_ (.D(_00277_),
    .CLK(clknet_leaf_173_clk),
    .Q(\channels.sample3[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17208_ (.D(_00278_),
    .CLK(clknet_5_24__leaf_clk),
    .Q(\channels.sample3[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17209_ (.D(_00279_),
    .CLK(clknet_leaf_94_clk),
    .Q(\channels.sample3[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17210_ (.D(_00280_),
    .CLK(clknet_leaf_93_clk),
    .Q(\channels.sample3[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17211_ (.D(_00281_),
    .CLK(clknet_leaf_94_clk),
    .Q(\channels.sample3[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17212_ (.D(_00282_),
    .CLK(clknet_leaf_171_clk),
    .Q(\channels.sample3[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17213_ (.D(_00283_),
    .CLK(clknet_leaf_170_clk),
    .Q(\channels.sample2[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17214_ (.D(_00284_),
    .CLK(clknet_leaf_179_clk),
    .Q(\channels.sample2[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17215_ (.D(_00285_),
    .CLK(clknet_leaf_179_clk),
    .Q(\channels.sample2[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17216_ (.D(_00286_),
    .CLK(clknet_leaf_175_clk),
    .Q(\channels.sample2[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17217_ (.D(_00287_),
    .CLK(clknet_leaf_174_clk),
    .Q(\channels.sample2[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17218_ (.D(_00288_),
    .CLK(clknet_leaf_174_clk),
    .Q(\channels.sample2[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17219_ (.D(_00289_),
    .CLK(clknet_leaf_173_clk),
    .Q(\channels.sample2[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17220_ (.D(_00290_),
    .CLK(clknet_leaf_173_clk),
    .Q(\channels.sample2[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17221_ (.D(_00291_),
    .CLK(clknet_leaf_94_clk),
    .Q(\channels.sample2[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17222_ (.D(_00292_),
    .CLK(clknet_leaf_93_clk),
    .Q(\channels.sample2[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17223_ (.D(_00293_),
    .CLK(clknet_leaf_93_clk),
    .Q(\channels.sample2[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17224_ (.D(_00294_),
    .CLK(clknet_leaf_169_clk),
    .Q(\channels.sample2[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17225_ (.D(_00295_),
    .CLK(clknet_leaf_170_clk),
    .Q(\channels.sample1[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17226_ (.D(_00296_),
    .CLK(clknet_leaf_176_clk),
    .Q(\channels.sample1[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17227_ (.D(_00297_),
    .CLK(clknet_leaf_176_clk),
    .Q(\channels.sample1[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17228_ (.D(_00298_),
    .CLK(clknet_leaf_176_clk),
    .Q(\channels.sample1[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17229_ (.D(_00299_),
    .CLK(clknet_leaf_174_clk),
    .Q(\channels.sample1[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17230_ (.D(_00300_),
    .CLK(clknet_leaf_173_clk),
    .Q(\channels.sample1[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17231_ (.D(_00301_),
    .CLK(clknet_leaf_170_clk),
    .Q(\channels.sample1[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17232_ (.D(_00302_),
    .CLK(clknet_leaf_172_clk),
    .Q(\channels.sample1[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17233_ (.D(_00303_),
    .CLK(clknet_leaf_172_clk),
    .Q(\channels.sample1[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17234_ (.D(_00304_),
    .CLK(clknet_leaf_171_clk),
    .Q(\channels.sample1[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17235_ (.D(_00305_),
    .CLK(clknet_leaf_171_clk),
    .Q(\channels.sample1[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17236_ (.D(_00306_),
    .CLK(clknet_leaf_170_clk),
    .Q(\channels.sample1[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17237_ (.D(_00307_),
    .CLK(clknet_5_6__leaf_clk),
    .Q(\filters.sample_filtered[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17238_ (.D(_00308_),
    .CLK(clknet_leaf_13_clk),
    .Q(\filters.sample_filtered[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17239_ (.D(_00309_),
    .CLK(clknet_leaf_91_clk),
    .Q(\filters.sample_filtered[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17240_ (.D(_00310_),
    .CLK(clknet_5_7__leaf_clk),
    .Q(\filters.sample_filtered[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17241_ (.D(_00311_),
    .CLK(clknet_leaf_11_clk),
    .Q(\filters.sample_filtered[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17242_ (.D(_00312_),
    .CLK(clknet_leaf_11_clk),
    .Q(\filters.sample_filtered[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17243_ (.D(_00313_),
    .CLK(clknet_leaf_91_clk),
    .Q(\filters.sample_filtered[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17244_ (.D(_00314_),
    .CLK(clknet_leaf_90_clk),
    .Q(\filters.sample_filtered[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17245_ (.D(_00315_),
    .CLK(clknet_leaf_90_clk),
    .Q(\filters.sample_filtered[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17246_ (.D(_00316_),
    .CLK(clknet_leaf_85_clk),
    .Q(\filters.sample_filtered[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17247_ (.D(_00317_),
    .CLK(clknet_leaf_86_clk),
    .Q(\filters.sample_filtered[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17248_ (.D(_00318_),
    .CLK(clknet_leaf_85_clk),
    .Q(\filters.sample_filtered[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17249_ (.D(_00319_),
    .CLK(clknet_leaf_91_clk),
    .Q(\filters.sample_filtered[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17250_ (.D(_00320_),
    .CLK(clknet_5_6__leaf_clk),
    .Q(\filters.sample_filtered[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17251_ (.D(_00321_),
    .CLK(clknet_leaf_86_clk),
    .Q(\filters.sample_filtered[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17252_ (.D(_00322_),
    .CLK(clknet_leaf_18_clk),
    .Q(\filters.sample_filtered[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17253_ (.D(_00323_),
    .CLK(clknet_leaf_75_clk),
    .Q(\filters.cutoff_lut[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17254_ (.D(_00324_),
    .CLK(clknet_leaf_75_clk),
    .Q(\filters.cutoff_lut[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17255_ (.D(_00325_),
    .CLK(clknet_leaf_76_clk),
    .Q(\filters.cutoff_lut[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17256_ (.D(_00326_),
    .CLK(clknet_leaf_73_clk),
    .Q(\tt_um_rejunity_sn76489.control_tone_freq[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17257_ (.D(_00327_),
    .CLK(clknet_leaf_71_clk),
    .Q(\tt_um_rejunity_sn76489.control_tone_freq[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17258_ (.D(_00328_),
    .CLK(clknet_leaf_72_clk),
    .Q(\tt_um_rejunity_sn76489.control_tone_freq[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17259_ (.D(_00329_),
    .CLK(clknet_leaf_72_clk),
    .Q(\tt_um_rejunity_sn76489.control_tone_freq[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17260_ (.D(_00330_),
    .CLK(clknet_leaf_74_clk),
    .Q(\tt_um_rejunity_sn76489.control_tone_freq[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17261_ (.D(_00331_),
    .CLK(clknet_leaf_75_clk),
    .Q(\tt_um_rejunity_sn76489.control_tone_freq[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17262_ (.D(_00332_),
    .CLK(clknet_leaf_75_clk),
    .Q(\tt_um_rejunity_sn76489.control_tone_freq[2][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17263_ (.D(_00333_),
    .CLK(clknet_leaf_75_clk),
    .Q(\tt_um_rejunity_sn76489.control_tone_freq[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17264_ (.D(_00334_),
    .CLK(clknet_leaf_71_clk),
    .Q(\tt_um_rejunity_sn76489.control_tone_freq[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17265_ (.D(_00335_),
    .CLK(clknet_leaf_70_clk),
    .Q(\tt_um_rejunity_sn76489.control_tone_freq[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17266_ (.D(_00336_),
    .CLK(clknet_leaf_70_clk),
    .Q(\tt_um_rejunity_sn76489.control_tone_freq[1][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17267_ (.D(_00337_),
    .CLK(clknet_leaf_70_clk),
    .Q(\tt_um_rejunity_sn76489.control_tone_freq[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17268_ (.D(_00338_),
    .CLK(clknet_leaf_153_clk),
    .Q(\channels.adsr_state[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17269_ (.D(_00339_),
    .CLK(clknet_leaf_153_clk),
    .Q(\channels.adsr_state[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17270_ (.D(_00340_),
    .CLK(clknet_leaf_182_clk),
    .Q(\channels.accum[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17271_ (.D(_00341_),
    .CLK(clknet_leaf_178_clk),
    .Q(\channels.accum[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17272_ (.D(_00342_),
    .CLK(clknet_leaf_187_clk),
    .Q(\channels.accum[2][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17273_ (.D(_00343_),
    .CLK(clknet_leaf_179_clk),
    .Q(\channels.accum[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17274_ (.D(_00344_),
    .CLK(clknet_leaf_186_clk),
    .Q(\channels.accum[2][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17275_ (.D(_00345_),
    .CLK(clknet_leaf_179_clk),
    .Q(\channels.accum[2][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17276_ (.D(_00346_),
    .CLK(clknet_leaf_181_clk),
    .Q(\channels.accum[2][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17277_ (.D(_00347_),
    .CLK(clknet_leaf_169_clk),
    .Q(\channels.accum[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17278_ (.D(_00348_),
    .CLK(clknet_leaf_153_clk),
    .Q(\channels.accum[2][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17279_ (.D(_00349_),
    .CLK(clknet_leaf_163_clk),
    .Q(\channels.accum[2][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17280_ (.D(_00350_),
    .CLK(clknet_leaf_147_clk),
    .Q(\channels.accum[2][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17281_ (.D(_00351_),
    .CLK(clknet_leaf_165_clk),
    .Q(\channels.accum[2][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17282_ (.D(_00352_),
    .CLK(clknet_leaf_152_clk),
    .Q(\channels.accum[2][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17283_ (.D(_00353_),
    .CLK(clknet_leaf_164_clk),
    .Q(\channels.accum[2][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17284_ (.D(_00354_),
    .CLK(clknet_leaf_154_clk),
    .Q(\channels.accum[2][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17285_ (.D(_00355_),
    .CLK(clknet_leaf_162_clk),
    .Q(\channels.accum[2][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17286_ (.D(_00356_),
    .CLK(clknet_leaf_158_clk),
    .Q(\channels.accum[2][16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17287_ (.D(_00357_),
    .CLK(clknet_leaf_190_clk),
    .Q(\channels.accum[2][17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17288_ (.D(_00358_),
    .CLK(clknet_leaf_157_clk),
    .Q(\channels.accum[2][18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17289_ (.D(_00359_),
    .CLK(clknet_leaf_161_clk),
    .Q(\channels.accum[2][19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17290_ (.D(_00360_),
    .CLK(clknet_leaf_158_clk),
    .Q(\channels.accum[2][20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17291_ (.D(_00361_),
    .CLK(clknet_leaf_189_clk),
    .Q(\channels.accum[2][21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17292_ (.D(_00362_),
    .CLK(clknet_leaf_155_clk),
    .Q(\channels.accum[2][22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17293_ (.D(_00363_),
    .CLK(clknet_leaf_188_clk),
    .Q(\channels.accum[2][23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17294_ (.D(_00364_),
    .CLK(clknet_leaf_187_clk),
    .Q(\channels.accum[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17295_ (.D(_00365_),
    .CLK(clknet_leaf_182_clk),
    .Q(\channels.accum[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17296_ (.D(_00366_),
    .CLK(clknet_leaf_186_clk),
    .Q(\channels.accum[1][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17297_ (.D(_00367_),
    .CLK(clknet_leaf_178_clk),
    .Q(\channels.accum[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17298_ (.D(_00368_),
    .CLK(clknet_leaf_186_clk),
    .Q(\channels.accum[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17299_ (.D(_00369_),
    .CLK(clknet_leaf_179_clk),
    .Q(\channels.accum[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17300_ (.D(_00370_),
    .CLK(clknet_leaf_188_clk),
    .Q(\channels.accum[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17301_ (.D(_00371_),
    .CLK(clknet_leaf_169_clk),
    .Q(\channels.accum[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17302_ (.D(_00372_),
    .CLK(clknet_leaf_154_clk),
    .Q(\channels.accum[1][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17303_ (.D(_00373_),
    .CLK(clknet_leaf_163_clk),
    .Q(\channels.accum[1][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17304_ (.D(_00374_),
    .CLK(clknet_leaf_152_clk),
    .Q(\channels.accum[1][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17305_ (.D(_00375_),
    .CLK(clknet_leaf_146_clk),
    .Q(\channels.accum[1][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17306_ (.D(_00376_),
    .CLK(clknet_leaf_152_clk),
    .Q(\channels.accum[1][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17307_ (.D(_00377_),
    .CLK(clknet_leaf_164_clk),
    .Q(\channels.accum[1][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17308_ (.D(_00378_),
    .CLK(clknet_leaf_154_clk),
    .Q(\channels.accum[1][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17309_ (.D(_00379_),
    .CLK(clknet_leaf_158_clk),
    .Q(\channels.accum[1][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17310_ (.D(_00380_),
    .CLK(clknet_leaf_156_clk),
    .Q(\channels.accum[1][16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17311_ (.D(_00381_),
    .CLK(clknet_leaf_192_clk),
    .Q(\channels.accum[1][17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17312_ (.D(_00382_),
    .CLK(clknet_leaf_157_clk),
    .Q(\channels.accum[1][18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17313_ (.D(_00383_),
    .CLK(clknet_leaf_161_clk),
    .Q(\channels.accum[1][19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17314_ (.D(_00384_),
    .CLK(clknet_leaf_157_clk),
    .Q(\channels.accum[1][20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17315_ (.D(_00385_),
    .CLK(clknet_leaf_190_clk),
    .Q(\channels.accum[1][21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17316_ (.D(_00386_),
    .CLK(clknet_leaf_156_clk),
    .Q(\channels.accum[1][22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17317_ (.D(_00387_),
    .CLK(clknet_leaf_189_clk),
    .Q(\channels.accum[1][23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17318_ (.D(_00388_),
    .CLK(clknet_leaf_243_clk),
    .Q(\filters.res_lut[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17319_ (.D(_00389_),
    .CLK(clknet_leaf_243_clk),
    .Q(\filters.res_lut[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17320_ (.D(_00390_),
    .CLK(clknet_leaf_77_clk),
    .Q(\channels.freq1[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17321_ (.D(_00391_),
    .CLK(clknet_leaf_87_clk),
    .Q(\channels.freq1[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17322_ (.D(_00392_),
    .CLK(clknet_leaf_77_clk),
    .Q(\channels.freq1[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17323_ (.D(_00393_),
    .CLK(clknet_leaf_77_clk),
    .Q(\channels.freq1[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17324_ (.D(_00394_),
    .CLK(clknet_leaf_88_clk),
    .Q(\channels.freq1[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17325_ (.D(_00395_),
    .CLK(clknet_leaf_99_clk),
    .Q(\channels.freq1[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17326_ (.D(_00396_),
    .CLK(clknet_leaf_87_clk),
    .Q(\channels.freq1[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17327_ (.D(_00397_),
    .CLK(clknet_leaf_88_clk),
    .Q(\channels.freq1[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17328_ (.D(_00398_),
    .CLK(clknet_leaf_87_clk),
    .Q(\channels.pw1[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17329_ (.D(_00399_),
    .CLK(clknet_leaf_87_clk),
    .Q(\channels.pw1[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17330_ (.D(_00400_),
    .CLK(clknet_leaf_86_clk),
    .Q(\channels.pw1[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17331_ (.D(_00401_),
    .CLK(clknet_leaf_86_clk),
    .Q(\channels.pw1[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17332_ (.D(_00402_),
    .CLK(clknet_leaf_97_clk),
    .Q(\channels.pw1[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17333_ (.D(_00403_),
    .CLK(clknet_leaf_89_clk),
    .Q(\channels.pw1[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17334_ (.D(_00404_),
    .CLK(clknet_leaf_89_clk),
    .Q(\channels.pw1[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17335_ (.D(_00405_),
    .CLK(clknet_leaf_97_clk),
    .Q(\channels.pw1[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17336_ (.D(_00406_),
    .CLK(clknet_leaf_100_clk),
    .Q(\channels.freq2[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17337_ (.D(_00407_),
    .CLK(clknet_leaf_103_clk),
    .Q(\channels.freq2[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17338_ (.D(_00408_),
    .CLK(clknet_leaf_103_clk),
    .Q(\channels.freq2[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17339_ (.D(_00409_),
    .CLK(clknet_leaf_103_clk),
    .Q(\channels.freq2[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17340_ (.D(_00410_),
    .CLK(clknet_leaf_100_clk),
    .Q(\channels.freq2[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17341_ (.D(_00411_),
    .CLK(clknet_leaf_102_clk),
    .Q(\channels.freq2[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17342_ (.D(_00412_),
    .CLK(clknet_leaf_100_clk),
    .Q(\channels.freq2[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17343_ (.D(_00413_),
    .CLK(clknet_leaf_102_clk),
    .Q(\channels.freq2[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17344_ (.D(_00414_),
    .CLK(clknet_leaf_100_clk),
    .Q(\channels.freq3[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17345_ (.D(_00415_),
    .CLK(clknet_leaf_96_clk),
    .Q(\channels.freq3[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17346_ (.D(_00416_),
    .CLK(clknet_leaf_98_clk),
    .Q(\channels.freq3[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17347_ (.D(_00417_),
    .CLK(clknet_leaf_100_clk),
    .Q(\channels.freq3[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17348_ (.D(_00418_),
    .CLK(clknet_leaf_101_clk),
    .Q(\channels.freq3[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17349_ (.D(_00419_),
    .CLK(clknet_leaf_100_clk),
    .Q(\channels.freq3[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17350_ (.D(_00420_),
    .CLK(clknet_leaf_101_clk),
    .Q(\channels.freq3[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17351_ (.D(_00421_),
    .CLK(clknet_leaf_101_clk),
    .Q(\channels.freq3[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17352_ (.D(_00422_),
    .CLK(clknet_leaf_96_clk),
    .Q(\channels.pw3[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17353_ (.D(_00423_),
    .CLK(clknet_leaf_96_clk),
    .Q(\channels.pw3[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17354_ (.D(_00424_),
    .CLK(clknet_leaf_96_clk),
    .Q(\channels.pw3[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17355_ (.D(_00425_),
    .CLK(clknet_leaf_95_clk),
    .Q(\channels.pw3[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17356_ (.D(_00426_),
    .CLK(clknet_leaf_172_clk),
    .Q(\channels.pw3[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17357_ (.D(_00427_),
    .CLK(clknet_leaf_101_clk),
    .Q(\channels.pw3[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17358_ (.D(_00428_),
    .CLK(clknet_leaf_95_clk),
    .Q(\channels.pw3[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17359_ (.D(_00429_),
    .CLK(clknet_leaf_172_clk),
    .Q(\channels.pw3[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17360_ (.D(_00430_),
    .CLK(clknet_leaf_89_clk),
    .Q(\channels.pw2[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17361_ (.D(_00431_),
    .CLK(clknet_leaf_97_clk),
    .Q(\channels.pw2[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17362_ (.D(_00432_),
    .CLK(clknet_leaf_93_clk),
    .Q(\channels.pw2[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17363_ (.D(_00433_),
    .CLK(clknet_leaf_97_clk),
    .Q(\channels.pw2[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17364_ (.D(_00434_),
    .CLK(clknet_leaf_171_clk),
    .Q(\channels.pw2[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17365_ (.D(_00435_),
    .CLK(clknet_5_25__leaf_clk),
    .Q(\channels.pw2[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17366_ (.D(_00436_),
    .CLK(clknet_leaf_101_clk),
    .Q(\channels.pw2[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17367_ (.D(_00437_),
    .CLK(clknet_leaf_171_clk),
    .Q(\channels.pw2[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _17368_ (.D(_00438_),
    .CLK(clknet_leaf_85_clk),
    .Q(\channels.clk_div[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17369_ (.D(_00439_),
    .CLK(clknet_leaf_165_clk),
    .Q(\channels.clk_div[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17370_ (.D(_00440_),
    .CLK(clknet_leaf_166_clk),
    .Q(\channels.clk_div[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17371_ (.D(_00441_),
    .CLK(clknet_leaf_209_clk),
    .Q(\channels.env_vol[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17372_ (.D(_00442_),
    .CLK(clknet_leaf_208_clk),
    .Q(\channels.env_vol[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17373_ (.D(_00443_),
    .CLK(clknet_leaf_210_clk),
    .Q(\channels.env_vol[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17374_ (.D(_00444_),
    .CLK(clknet_leaf_207_clk),
    .Q(\channels.env_vol[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17375_ (.D(_00445_),
    .CLK(clknet_leaf_204_clk),
    .Q(\channels.env_vol[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17376_ (.D(_00446_),
    .CLK(clknet_leaf_207_clk),
    .Q(\channels.env_vol[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17377_ (.D(_00447_),
    .CLK(clknet_leaf_214_clk),
    .Q(\channels.env_vol[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17378_ (.D(_00448_),
    .CLK(clknet_leaf_204_clk),
    .Q(\channels.env_vol[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17379_ (.D(_00449_),
    .CLK(clknet_leaf_131_clk),
    .Q(\channels.env_counter[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17380_ (.D(_00450_),
    .CLK(clknet_leaf_132_clk),
    .Q(\channels.env_counter[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17381_ (.D(_00451_),
    .CLK(clknet_leaf_134_clk),
    .Q(\channels.env_counter[2][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17382_ (.D(_00452_),
    .CLK(clknet_leaf_129_clk),
    .Q(\channels.env_counter[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17383_ (.D(_00453_),
    .CLK(clknet_leaf_136_clk),
    .Q(\channels.env_counter[2][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17384_ (.D(_00454_),
    .CLK(clknet_leaf_137_clk),
    .Q(\channels.env_counter[2][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17385_ (.D(_00455_),
    .CLK(clknet_5_31__leaf_clk),
    .Q(\channels.env_counter[2][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17386_ (.D(_00456_),
    .CLK(clknet_leaf_136_clk),
    .Q(\channels.env_counter[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17387_ (.D(_00457_),
    .CLK(clknet_leaf_149_clk),
    .Q(\channels.env_counter[2][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17388_ (.D(_00458_),
    .CLK(clknet_leaf_149_clk),
    .Q(\channels.env_counter[2][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17389_ (.D(_00459_),
    .CLK(clknet_leaf_148_clk),
    .Q(\channels.env_counter[2][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17390_ (.D(_00460_),
    .CLK(clknet_leaf_148_clk),
    .Q(\channels.env_counter[2][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17391_ (.D(_00461_),
    .CLK(clknet_leaf_123_clk),
    .Q(\channels.env_counter[2][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17392_ (.D(_00462_),
    .CLK(clknet_leaf_130_clk),
    .Q(\channels.env_counter[2][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17393_ (.D(_00463_),
    .CLK(clknet_leaf_129_clk),
    .Q(\channels.env_counter[2][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17394_ (.D(_00464_),
    .CLK(clknet_leaf_132_clk),
    .Q(\channels.env_counter[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17395_ (.D(_00465_),
    .CLK(clknet_leaf_132_clk),
    .Q(\channels.env_counter[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17396_ (.D(_00466_),
    .CLK(clknet_leaf_132_clk),
    .Q(\channels.env_counter[1][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17397_ (.D(_00467_),
    .CLK(clknet_leaf_131_clk),
    .Q(\channels.env_counter[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17398_ (.D(_00468_),
    .CLK(clknet_leaf_135_clk),
    .Q(\channels.env_counter[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17399_ (.D(_00469_),
    .CLK(clknet_leaf_138_clk),
    .Q(\channels.env_counter[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17400_ (.D(_00470_),
    .CLK(clknet_leaf_139_clk),
    .Q(\channels.env_counter[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17401_ (.D(_00471_),
    .CLK(clknet_leaf_137_clk),
    .Q(\channels.env_counter[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17402_ (.D(_00472_),
    .CLK(clknet_leaf_150_clk),
    .Q(\channels.env_counter[1][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17403_ (.D(_00473_),
    .CLK(clknet_leaf_149_clk),
    .Q(\channels.env_counter[1][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17404_ (.D(_00474_),
    .CLK(clknet_leaf_148_clk),
    .Q(\channels.env_counter[1][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17405_ (.D(_00475_),
    .CLK(clknet_leaf_149_clk),
    .Q(\channels.env_counter[1][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17406_ (.D(_00476_),
    .CLK(clknet_leaf_130_clk),
    .Q(\channels.env_counter[1][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17407_ (.D(_00477_),
    .CLK(clknet_leaf_130_clk),
    .Q(\channels.env_counter[1][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17408_ (.D(_00478_),
    .CLK(clknet_leaf_129_clk),
    .Q(\channels.env_counter[1][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17409_ (.D(_00479_),
    .CLK(clknet_leaf_158_clk),
    .Q(\channels.adsr_state[3][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17410_ (.D(_00480_),
    .CLK(clknet_leaf_147_clk),
    .Q(\channels.adsr_state[3][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17411_ (.D(_00481_),
    .CLK(clknet_leaf_86_clk),
    .Q(\clk_ctr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17412_ (.D(_00482_),
    .CLK(clknet_leaf_86_clk),
    .Q(\clk_ctr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17413_ (.D(_00483_),
    .CLK(clknet_leaf_132_clk),
    .Q(\channels.env_counter[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17414_ (.D(_00484_),
    .CLK(clknet_leaf_132_clk),
    .Q(\channels.env_counter[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17415_ (.D(_00485_),
    .CLK(clknet_leaf_134_clk),
    .Q(\channels.env_counter[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17416_ (.D(_00486_),
    .CLK(clknet_leaf_131_clk),
    .Q(\channels.env_counter[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17417_ (.D(_00487_),
    .CLK(clknet_leaf_135_clk),
    .Q(\channels.env_counter[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17418_ (.D(_00488_),
    .CLK(clknet_leaf_138_clk),
    .Q(\channels.env_counter[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17419_ (.D(_00489_),
    .CLK(clknet_leaf_139_clk),
    .Q(\channels.env_counter[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17420_ (.D(_00490_),
    .CLK(clknet_leaf_137_clk),
    .Q(\channels.env_counter[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17421_ (.D(_00491_),
    .CLK(clknet_leaf_150_clk),
    .Q(\channels.env_counter[0][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17422_ (.D(_00492_),
    .CLK(clknet_leaf_150_clk),
    .Q(\channels.env_counter[0][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17423_ (.D(_00493_),
    .CLK(clknet_leaf_149_clk),
    .Q(\channels.env_counter[0][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17424_ (.D(_00494_),
    .CLK(clknet_leaf_148_clk),
    .Q(\channels.env_counter[0][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17425_ (.D(_00495_),
    .CLK(clknet_leaf_130_clk),
    .Q(\channels.env_counter[0][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17426_ (.D(_00496_),
    .CLK(clknet_leaf_136_clk),
    .Q(\channels.env_counter[0][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17427_ (.D(_00497_),
    .CLK(clknet_leaf_129_clk),
    .Q(\channels.env_counter[0][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17428_ (.D(_00498_),
    .CLK(clknet_leaf_159_clk),
    .Q(\channels.adsr_state[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17429_ (.D(_00499_),
    .CLK(clknet_leaf_164_clk),
    .Q(\channels.adsr_state[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17430_ (.D(_00500_),
    .CLK(clknet_leaf_159_clk),
    .Q(\channels.adsr_state[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17431_ (.D(_00501_),
    .CLK(clknet_leaf_153_clk),
    .Q(\channels.adsr_state[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17432_ (.D(_00502_),
    .CLK(clknet_leaf_182_clk),
    .Q(\channels.accum[3][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17433_ (.D(_00503_),
    .CLK(clknet_leaf_182_clk),
    .Q(\channels.accum[3][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17434_ (.D(_00504_),
    .CLK(clknet_leaf_187_clk),
    .Q(\channels.accum[3][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17435_ (.D(_00505_),
    .CLK(clknet_leaf_178_clk),
    .Q(\channels.accum[3][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17436_ (.D(_00506_),
    .CLK(clknet_leaf_185_clk),
    .Q(\channels.accum[3][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17437_ (.D(_00507_),
    .CLK(clknet_leaf_180_clk),
    .Q(\channels.accum[3][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17438_ (.D(_00508_),
    .CLK(clknet_leaf_181_clk),
    .Q(\channels.accum[3][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17439_ (.D(_00509_),
    .CLK(clknet_leaf_169_clk),
    .Q(\channels.accum[3][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17440_ (.D(_00510_),
    .CLK(clknet_leaf_153_clk),
    .Q(\channels.accum[3][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17441_ (.D(_00511_),
    .CLK(clknet_leaf_163_clk),
    .Q(\channels.accum[3][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17442_ (.D(_00512_),
    .CLK(clknet_leaf_147_clk),
    .Q(\channels.accum[3][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17443_ (.D(_00513_),
    .CLK(clknet_leaf_146_clk),
    .Q(\channels.accum[3][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17444_ (.D(_00514_),
    .CLK(clknet_leaf_151_clk),
    .Q(\channels.accum[3][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17445_ (.D(_00515_),
    .CLK(clknet_leaf_147_clk),
    .Q(\channels.accum[3][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17446_ (.D(_00516_),
    .CLK(clknet_leaf_151_clk),
    .Q(\channels.accum[3][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17447_ (.D(_00517_),
    .CLK(clknet_leaf_162_clk),
    .Q(\channels.accum[3][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17448_ (.D(_00518_),
    .CLK(clknet_leaf_158_clk),
    .Q(\channels.accum[3][16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17449_ (.D(_00519_),
    .CLK(clknet_leaf_190_clk),
    .Q(\channels.accum[3][17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17450_ (.D(_00520_),
    .CLK(clknet_leaf_195_clk),
    .Q(\channels.accum[3][18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17451_ (.D(_00521_),
    .CLK(clknet_leaf_158_clk),
    .Q(\channels.accum[3][19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17452_ (.D(_00522_),
    .CLK(clknet_leaf_157_clk),
    .Q(\channels.accum[3][20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17453_ (.D(_00523_),
    .CLK(clknet_leaf_191_clk),
    .Q(\channels.accum[3][21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17454_ (.D(_00524_),
    .CLK(clknet_leaf_155_clk),
    .Q(\channels.accum[3][22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17455_ (.D(_00525_),
    .CLK(clknet_leaf_188_clk),
    .Q(\channels.accum[3][23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17456_ (.D(_00526_),
    .CLK(clknet_leaf_0_clk),
    .Q(\filters.band[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17457_ (.D(_00527_),
    .CLK(clknet_leaf_4_clk),
    .Q(\filters.band[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17458_ (.D(_00528_),
    .CLK(clknet_leaf_1_clk),
    .Q(\filters.band[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17459_ (.D(_00529_),
    .CLK(clknet_leaf_4_clk),
    .Q(\filters.band[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17460_ (.D(_00530_),
    .CLK(clknet_leaf_249_clk),
    .Q(\filters.band[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17461_ (.D(_00531_),
    .CLK(clknet_leaf_1_clk),
    .Q(\filters.band[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17462_ (.D(_00532_),
    .CLK(clknet_leaf_2_clk),
    .Q(\filters.band[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17463_ (.D(_00533_),
    .CLK(clknet_leaf_1_clk),
    .Q(\filters.band[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17464_ (.D(_00534_),
    .CLK(clknet_leaf_2_clk),
    .Q(\filters.band[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17465_ (.D(_00535_),
    .CLK(clknet_leaf_2_clk),
    .Q(\filters.band[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17466_ (.D(_00536_),
    .CLK(clknet_5_1__leaf_clk),
    .Q(\filters.band[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17467_ (.D(_00537_),
    .CLK(clknet_leaf_26_clk),
    .Q(\filters.band[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17468_ (.D(_00538_),
    .CLK(clknet_leaf_26_clk),
    .Q(\filters.band[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17469_ (.D(_00539_),
    .CLK(clknet_leaf_15_clk),
    .Q(\filters.band[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17470_ (.D(_00540_),
    .CLK(clknet_leaf_15_clk),
    .Q(\filters.band[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17471_ (.D(_00541_),
    .CLK(clknet_leaf_21_clk),
    .Q(\filters.band[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17472_ (.D(_00542_),
    .CLK(clknet_leaf_245_clk),
    .Q(\filters.band[16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17473_ (.D(_00543_),
    .CLK(clknet_leaf_27_clk),
    .Q(\filters.band[17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17474_ (.D(_00544_),
    .CLK(clknet_leaf_244_clk),
    .Q(\filters.band[18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17475_ (.D(_00545_),
    .CLK(clknet_leaf_244_clk),
    .Q(\filters.band[19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17476_ (.D(_00546_),
    .CLK(clknet_leaf_245_clk),
    .Q(\filters.band[20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17477_ (.D(_00547_),
    .CLK(clknet_leaf_29_clk),
    .Q(\filters.band[21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17478_ (.D(_00548_),
    .CLK(clknet_leaf_29_clk),
    .Q(\filters.band[22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17479_ (.D(_00549_),
    .CLK(clknet_leaf_29_clk),
    .Q(\filters.band[23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17480_ (.D(_00550_),
    .CLK(clknet_leaf_23_clk),
    .Q(\filters.band[24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17481_ (.D(_00551_),
    .CLK(clknet_leaf_32_clk),
    .Q(\filters.band[25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17482_ (.D(_00552_),
    .CLK(clknet_leaf_244_clk),
    .Q(\filters.band[26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17483_ (.D(_00553_),
    .CLK(clknet_leaf_244_clk),
    .Q(\filters.band[27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17484_ (.D(_00554_),
    .CLK(clknet_leaf_244_clk),
    .Q(\filters.band[28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17485_ (.D(_00555_),
    .CLK(clknet_leaf_246_clk),
    .Q(\filters.band[29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17486_ (.D(_00556_),
    .CLK(clknet_leaf_27_clk),
    .Q(\filters.band[30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17487_ (.D(_00557_),
    .CLK(clknet_leaf_23_clk),
    .Q(\filters.band[31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17488_ (.D(_00558_),
    .CLK(clknet_leaf_13_clk),
    .Q(\filters.high[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17489_ (.D(_00559_),
    .CLK(clknet_leaf_13_clk),
    .Q(\filters.high[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17490_ (.D(_00560_),
    .CLK(clknet_leaf_13_clk),
    .Q(\filters.high[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17491_ (.D(_00561_),
    .CLK(clknet_leaf_243_clk),
    .Q(\filters.high[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17492_ (.D(_00562_),
    .CLK(clknet_leaf_8_clk),
    .Q(\filters.high[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17493_ (.D(_00563_),
    .CLK(clknet_leaf_6_clk),
    .Q(\filters.high[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17494_ (.D(_00564_),
    .CLK(clknet_leaf_249_clk),
    .Q(\filters.high[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17495_ (.D(_00565_),
    .CLK(clknet_5_5__leaf_clk),
    .Q(\filters.high[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17496_ (.D(_00566_),
    .CLK(clknet_leaf_9_clk),
    .Q(\filters.high[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17497_ (.D(_00567_),
    .CLK(clknet_leaf_9_clk),
    .Q(\filters.high[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17498_ (.D(_00568_),
    .CLK(clknet_leaf_13_clk),
    .Q(\filters.high[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17499_ (.D(_00569_),
    .CLK(clknet_leaf_6_clk),
    .Q(\filters.high[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17500_ (.D(_00570_),
    .CLK(clknet_leaf_249_clk),
    .Q(\filters.high[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17501_ (.D(_00571_),
    .CLK(clknet_leaf_14_clk),
    .Q(\filters.high[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17502_ (.D(_00572_),
    .CLK(clknet_leaf_14_clk),
    .Q(\filters.high[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17503_ (.D(_00573_),
    .CLK(clknet_leaf_21_clk),
    .Q(\filters.high[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17504_ (.D(_00574_),
    .CLK(clknet_leaf_248_clk),
    .Q(\filters.high[16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17505_ (.D(_00575_),
    .CLK(clknet_leaf_249_clk),
    .Q(\filters.high[17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17506_ (.D(_00576_),
    .CLK(clknet_leaf_248_clk),
    .Q(\filters.high[18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17507_ (.D(_00577_),
    .CLK(clknet_leaf_247_clk),
    .Q(\filters.high[19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17508_ (.D(_00578_),
    .CLK(clknet_leaf_247_clk),
    .Q(\filters.high[20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17509_ (.D(_00579_),
    .CLK(clknet_leaf_246_clk),
    .Q(\filters.high[21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17510_ (.D(_00580_),
    .CLK(clknet_leaf_27_clk),
    .Q(\filters.high[22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17511_ (.D(_00581_),
    .CLK(clknet_leaf_27_clk),
    .Q(\filters.high[23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17512_ (.D(_00582_),
    .CLK(clknet_leaf_27_clk),
    .Q(\filters.high[24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17513_ (.D(_00583_),
    .CLK(clknet_leaf_21_clk),
    .Q(\filters.high[25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17514_ (.D(_00584_),
    .CLK(clknet_leaf_21_clk),
    .Q(\filters.high[26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17515_ (.D(_00585_),
    .CLK(clknet_leaf_37_clk),
    .Q(\filters.high[27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17516_ (.D(_00586_),
    .CLK(clknet_5_1__leaf_clk),
    .Q(\filters.high[28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17517_ (.D(_00587_),
    .CLK(clknet_5_2__leaf_clk),
    .Q(\filters.high[29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17518_ (.D(_00588_),
    .CLK(clknet_leaf_37_clk),
    .Q(\filters.high[30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17519_ (.D(_00589_),
    .CLK(clknet_leaf_22_clk),
    .Q(\filters.high[31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17520_ (.D(_00590_),
    .CLK(clknet_leaf_18_clk),
    .Q(\filters.sample_buff[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17521_ (.D(_00591_),
    .CLK(clknet_leaf_18_clk),
    .Q(\filters.sample_buff[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17522_ (.D(_00592_),
    .CLK(clknet_leaf_21_clk),
    .Q(\filters.sample_buff[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17523_ (.D(_00593_),
    .CLK(clknet_leaf_20_clk),
    .Q(\filters.sample_buff[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17524_ (.D(_00594_),
    .CLK(clknet_leaf_19_clk),
    .Q(\filters.sample_buff[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17525_ (.D(_00595_),
    .CLK(clknet_leaf_20_clk),
    .Q(\filters.sample_buff[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17526_ (.D(_00596_),
    .CLK(clknet_leaf_19_clk),
    .Q(\filters.sample_buff[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17527_ (.D(_00597_),
    .CLK(clknet_leaf_19_clk),
    .Q(\filters.sample_buff[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17528_ (.D(_00598_),
    .CLK(clknet_5_6__leaf_clk),
    .Q(\filters.sample_buff[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17529_ (.D(_00599_),
    .CLK(clknet_leaf_82_clk),
    .Q(\filters.sample_buff[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17530_ (.D(_00600_),
    .CLK(clknet_leaf_82_clk),
    .Q(\filters.sample_buff[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17531_ (.D(_00601_),
    .CLK(clknet_leaf_82_clk),
    .Q(\filters.sample_buff[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17532_ (.D(_00602_),
    .CLK(clknet_leaf_82_clk),
    .Q(\filters.sample_buff[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17533_ (.D(_00603_),
    .CLK(clknet_leaf_82_clk),
    .Q(\filters.sample_buff[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17534_ (.D(_00604_),
    .CLK(clknet_leaf_20_clk),
    .Q(\filters.sample_buff[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17535_ (.D(_00605_),
    .CLK(clknet_leaf_200_clk),
    .Q(\channels.exp_periods[3][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17536_ (.D(_00606_),
    .CLK(clknet_leaf_215_clk),
    .Q(\channels.exp_periods[3][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17537_ (.D(_00607_),
    .CLK(clknet_leaf_215_clk),
    .Q(\channels.exp_periods[3][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17538_ (.D(_00608_),
    .CLK(clknet_leaf_202_clk),
    .Q(\channels.exp_periods[3][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17539_ (.D(_00609_),
    .CLK(clknet_leaf_201_clk),
    .Q(\channels.exp_periods[3][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17540_ (.D(_00610_),
    .CLK(clknet_leaf_5_clk),
    .Q(\filters.low[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17541_ (.D(_00611_),
    .CLK(clknet_leaf_5_clk),
    .Q(\filters.low[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17542_ (.D(_00612_),
    .CLK(clknet_leaf_243_clk),
    .Q(\filters.low[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17543_ (.D(_00613_),
    .CLK(clknet_leaf_243_clk),
    .Q(\filters.low[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17544_ (.D(_00614_),
    .CLK(clknet_leaf_0_clk),
    .Q(\filters.low[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17545_ (.D(_00615_),
    .CLK(clknet_leaf_242_clk),
    .Q(\filters.low[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17546_ (.D(_00616_),
    .CLK(clknet_leaf_242_clk),
    .Q(\filters.low[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17547_ (.D(_00617_),
    .CLK(clknet_leaf_242_clk),
    .Q(\filters.low[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17548_ (.D(_00618_),
    .CLK(clknet_leaf_8_clk),
    .Q(\filters.low[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17549_ (.D(_00619_),
    .CLK(clknet_leaf_175_clk),
    .Q(\filters.low[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17550_ (.D(_00620_),
    .CLK(clknet_leaf_5_clk),
    .Q(\filters.low[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17551_ (.D(_00621_),
    .CLK(clknet_leaf_14_clk),
    .Q(\filters.low[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17552_ (.D(_00622_),
    .CLK(clknet_leaf_14_clk),
    .Q(\filters.low[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17553_ (.D(_00623_),
    .CLK(clknet_leaf_25_clk),
    .Q(\filters.low[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17554_ (.D(_00624_),
    .CLK(clknet_leaf_25_clk),
    .Q(\filters.low[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17555_ (.D(_00625_),
    .CLK(clknet_leaf_23_clk),
    .Q(\filters.low[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17556_ (.D(_00626_),
    .CLK(clknet_leaf_246_clk),
    .Q(\filters.low[16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17557_ (.D(_00627_),
    .CLK(clknet_leaf_27_clk),
    .Q(\filters.low[17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17558_ (.D(_00628_),
    .CLK(clknet_leaf_244_clk),
    .Q(\filters.low[18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17559_ (.D(_00629_),
    .CLK(clknet_leaf_245_clk),
    .Q(\filters.low[19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17560_ (.D(_00630_),
    .CLK(clknet_leaf_29_clk),
    .Q(\filters.low[20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17561_ (.D(_00631_),
    .CLK(clknet_leaf_30_clk),
    .Q(\filters.low[21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17562_ (.D(_00632_),
    .CLK(clknet_leaf_30_clk),
    .Q(\filters.low[22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17563_ (.D(_00633_),
    .CLK(clknet_5_0__leaf_clk),
    .Q(\filters.low[23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17564_ (.D(_00634_),
    .CLK(clknet_5_2__leaf_clk),
    .Q(\filters.low[24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17565_ (.D(_00635_),
    .CLK(clknet_leaf_32_clk),
    .Q(\filters.low[25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17566_ (.D(_00636_),
    .CLK(clknet_leaf_32_clk),
    .Q(\filters.low[26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17567_ (.D(_00637_),
    .CLK(clknet_leaf_32_clk),
    .Q(\filters.low[27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17568_ (.D(_00638_),
    .CLK(clknet_leaf_34_clk),
    .Q(\filters.low[28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17569_ (.D(_00639_),
    .CLK(clknet_leaf_34_clk),
    .Q(\filters.low[29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17570_ (.D(_00640_),
    .CLK(clknet_leaf_37_clk),
    .Q(\filters.low[30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17571_ (.D(_00641_),
    .CLK(clknet_leaf_22_clk),
    .Q(\filters.low[31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17572_ (.D(_00642_),
    .CLK(clknet_5_5__leaf_clk),
    .Q(\filters.filter_step[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _17573_ (.D(_00643_),
    .CLK(clknet_5_5__leaf_clk),
    .Q(\filters.filter_step[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _17574_ (.D(_00644_),
    .CLK(clknet_leaf_6_clk),
    .Q(\filters.filter_step[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17575_ (.D(_00645_),
    .CLK(clknet_leaf_38_clk),
    .Q(\spi_dac_i.counter[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17576_ (.D(_00646_),
    .CLK(clknet_leaf_33_clk),
    .Q(\spi_dac_i.counter[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17577_ (.D(_00647_),
    .CLK(clknet_leaf_33_clk),
    .Q(\spi_dac_i.counter[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17578_ (.D(_00648_),
    .CLK(clknet_leaf_34_clk),
    .Q(\spi_dac_i.counter[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17579_ (.D(_00649_),
    .CLK(clknet_leaf_34_clk),
    .Q(\spi_dac_i.counter[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17580_ (.D(_00650_),
    .CLK(clknet_leaf_44_clk),
    .Q(\spi_dac_i.spi_dat_buff_1[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17581_ (.D(_00651_),
    .CLK(clknet_leaf_45_clk),
    .Q(\spi_dac_i.spi_dat_buff_1[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17582_ (.D(_00652_),
    .CLK(clknet_leaf_46_clk),
    .Q(\spi_dac_i.spi_dat_buff_1[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17583_ (.D(_00653_),
    .CLK(clknet_leaf_33_clk),
    .Q(\spi_dac_i.spi_dat_buff_1[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17584_ (.D(_00654_),
    .CLK(clknet_leaf_46_clk),
    .Q(\spi_dac_i.spi_dat_buff_1[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17585_ (.D(_00655_),
    .CLK(clknet_leaf_46_clk),
    .Q(\spi_dac_i.spi_dat_buff_1[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17586_ (.D(_00656_),
    .CLK(clknet_leaf_45_clk),
    .Q(\spi_dac_i.spi_dat_buff_1[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17587_ (.D(_00657_),
    .CLK(clknet_leaf_45_clk),
    .Q(\spi_dac_i.spi_dat_buff_1[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17588_ (.D(_00658_),
    .CLK(clknet_leaf_44_clk),
    .Q(\spi_dac_i.spi_dat_buff_1[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17589_ (.D(_00659_),
    .CLK(clknet_leaf_44_clk),
    .Q(\spi_dac_i.spi_dat_buff_1[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17590_ (.D(_00660_),
    .CLK(clknet_leaf_42_clk),
    .Q(\spi_dac_i.spi_dat_buff_1[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17591_ (.D(_00661_),
    .CLK(clknet_leaf_42_clk),
    .Q(\spi_dac_i.spi_dat_buff_1[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17592_ (.D(_00662_),
    .CLK(clknet_leaf_38_clk),
    .Q(\spi_dac_i.spi_dat_buff_0[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17593_ (.D(_00663_),
    .CLK(clknet_leaf_38_clk),
    .Q(\spi_dac_i.spi_dat_buff_0[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17594_ (.D(_00664_),
    .CLK(clknet_leaf_39_clk),
    .Q(\spi_dac_i.spi_dat_buff_0[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17595_ (.D(_00665_),
    .CLK(clknet_leaf_39_clk),
    .Q(\spi_dac_i.spi_dat_buff_0[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17596_ (.D(_00666_),
    .CLK(clknet_leaf_39_clk),
    .Q(\spi_dac_i.spi_dat_buff_0[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17597_ (.D(_00667_),
    .CLK(clknet_leaf_40_clk),
    .Q(\spi_dac_i.spi_dat_buff_0[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17598_ (.D(_00668_),
    .CLK(clknet_leaf_58_clk),
    .Q(\spi_dac_i.spi_dat_buff_0[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17599_ (.D(_00669_),
    .CLK(clknet_leaf_57_clk),
    .Q(\spi_dac_i.spi_dat_buff_0[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17600_ (.D(_00670_),
    .CLK(clknet_leaf_40_clk),
    .Q(\spi_dac_i.spi_dat_buff_0[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17601_ (.D(_00671_),
    .CLK(clknet_leaf_41_clk),
    .Q(\spi_dac_i.spi_dat_buff_0[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17602_ (.D(_00672_),
    .CLK(clknet_leaf_41_clk),
    .Q(\spi_dac_i.spi_dat_buff_0[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17603_ (.D(_00673_),
    .CLK(clknet_leaf_41_clk),
    .Q(\spi_dac_i.spi_dat_buff_0[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17604_ (.D(_00674_),
    .CLK(clknet_leaf_44_clk),
    .Q(net20));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17605_ (.D(_00675_),
    .CLK(clknet_leaf_44_clk),
    .Q(net19));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17606_ (.D(_00676_),
    .CLK(clknet_leaf_48_clk),
    .Q(net21));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17607_ (.D(_00677_),
    .CLK(clknet_leaf_162_clk),
    .Q(_00009_));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17608_ (.D(_00678_),
    .CLK(clknet_leaf_168_clk),
    .Q(_00010_));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17609_ (.D(_00679_),
    .CLK(clknet_leaf_131_clk),
    .Q(\channels.env_counter[3][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17610_ (.D(_00680_),
    .CLK(clknet_leaf_133_clk),
    .Q(\channels.env_counter[3][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17611_ (.D(_00681_),
    .CLK(clknet_leaf_133_clk),
    .Q(\channels.env_counter[3][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17612_ (.D(_00682_),
    .CLK(clknet_leaf_129_clk),
    .Q(\channels.env_counter[3][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17613_ (.D(_00683_),
    .CLK(clknet_leaf_135_clk),
    .Q(\channels.env_counter[3][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17614_ (.D(_00684_),
    .CLK(clknet_leaf_139_clk),
    .Q(\channels.env_counter[3][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17615_ (.D(_00685_),
    .CLK(clknet_leaf_139_clk),
    .Q(\channels.env_counter[3][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17616_ (.D(_00686_),
    .CLK(clknet_leaf_138_clk),
    .Q(\channels.env_counter[3][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17617_ (.D(_00687_),
    .CLK(clknet_leaf_150_clk),
    .Q(\channels.env_counter[3][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17618_ (.D(_00688_),
    .CLK(clknet_leaf_139_clk),
    .Q(\channels.env_counter[3][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17619_ (.D(_00689_),
    .CLK(clknet_leaf_145_clk),
    .Q(\channels.env_counter[3][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17620_ (.D(_00690_),
    .CLK(clknet_leaf_147_clk),
    .Q(\channels.env_counter[3][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17621_ (.D(_00691_),
    .CLK(clknet_leaf_128_clk),
    .Q(\channels.env_counter[3][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17622_ (.D(_00692_),
    .CLK(clknet_leaf_133_clk),
    .Q(\channels.env_counter[3][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17623_ (.D(_00693_),
    .CLK(clknet_leaf_128_clk),
    .Q(\channels.env_counter[3][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17624_ (.D(_00694_),
    .CLK(clknet_leaf_209_clk),
    .Q(\channels.env_vol[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17625_ (.D(_00695_),
    .CLK(clknet_leaf_209_clk),
    .Q(\channels.env_vol[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17626_ (.D(_00696_),
    .CLK(clknet_leaf_209_clk),
    .Q(\channels.env_vol[1][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17627_ (.D(_00697_),
    .CLK(clknet_leaf_208_clk),
    .Q(\channels.env_vol[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17628_ (.D(_00698_),
    .CLK(clknet_leaf_213_clk),
    .Q(\channels.env_vol[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17629_ (.D(_00699_),
    .CLK(clknet_leaf_210_clk),
    .Q(\channels.env_vol[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17630_ (.D(_00700_),
    .CLK(clknet_leaf_213_clk),
    .Q(\channels.env_vol[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17631_ (.D(_00701_),
    .CLK(clknet_leaf_204_clk),
    .Q(\channels.env_vol[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17632_ (.D(_00702_),
    .CLK(clknet_leaf_195_clk),
    .Q(\channels.exp_counter[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17633_ (.D(_00703_),
    .CLK(clknet_leaf_195_clk),
    .Q(\channels.exp_counter[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17634_ (.D(_00704_),
    .CLK(clknet_leaf_197_clk),
    .Q(\channels.exp_counter[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17635_ (.D(_00705_),
    .CLK(clknet_5_23__leaf_clk),
    .Q(\channels.exp_counter[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17636_ (.D(_00706_),
    .CLK(clknet_leaf_185_clk),
    .Q(\channels.exp_counter[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17637_ (.D(_00707_),
    .CLK(clknet_leaf_208_clk),
    .Q(\channels.ch3_env[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17638_ (.D(_00708_),
    .CLK(clknet_5_19__leaf_clk),
    .Q(\channels.ch3_env[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17639_ (.D(_00709_),
    .CLK(clknet_leaf_208_clk),
    .Q(\channels.ch3_env[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17640_ (.D(_00710_),
    .CLK(clknet_leaf_207_clk),
    .Q(\channels.ch3_env[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17641_ (.D(_00711_),
    .CLK(clknet_leaf_204_clk),
    .Q(\channels.ch3_env[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17642_ (.D(_00712_),
    .CLK(clknet_leaf_206_clk),
    .Q(\channels.ch3_env[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17643_ (.D(_00713_),
    .CLK(clknet_leaf_206_clk),
    .Q(\channels.ch3_env[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17644_ (.D(_00714_),
    .CLK(clknet_leaf_206_clk),
    .Q(\channels.ch3_env[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17645_ (.D(_00715_),
    .CLK(clknet_leaf_49_clk),
    .Q(\tt_um_rejunity_sn76489.chan[3].attenuation.in ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17646_ (.D(_00716_),
    .CLK(clknet_leaf_51_clk),
    .Q(\tt_um_rejunity_sn76489.noise[0].gen.lfsr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17647_ (.D(_00717_),
    .CLK(clknet_leaf_50_clk),
    .Q(\tt_um_rejunity_sn76489.noise[0].gen.lfsr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17648_ (.D(_00718_),
    .CLK(clknet_leaf_50_clk),
    .Q(\tt_um_rejunity_sn76489.noise[0].gen.lfsr[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17649_ (.D(_00719_),
    .CLK(clknet_leaf_50_clk),
    .Q(\tt_um_rejunity_sn76489.noise[0].gen.lfsr[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17650_ (.D(_00720_),
    .CLK(clknet_leaf_51_clk),
    .Q(\tt_um_rejunity_sn76489.noise[0].gen.lfsr[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17651_ (.D(_00721_),
    .CLK(clknet_leaf_51_clk),
    .Q(\tt_um_rejunity_sn76489.noise[0].gen.lfsr[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17652_ (.D(_00722_),
    .CLK(clknet_leaf_51_clk),
    .Q(\tt_um_rejunity_sn76489.noise[0].gen.lfsr[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17653_ (.D(_00723_),
    .CLK(clknet_leaf_51_clk),
    .Q(\tt_um_rejunity_sn76489.noise[0].gen.lfsr[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17654_ (.D(_00724_),
    .CLK(clknet_leaf_64_clk),
    .Q(\tt_um_rejunity_sn76489.noise[0].gen.lfsr[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17655_ (.D(_00725_),
    .CLK(clknet_leaf_52_clk),
    .Q(\tt_um_rejunity_sn76489.noise[0].gen.lfsr[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17656_ (.D(_00726_),
    .CLK(clknet_leaf_52_clk),
    .Q(\tt_um_rejunity_sn76489.noise[0].gen.lfsr[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17657_ (.D(_00727_),
    .CLK(clknet_leaf_52_clk),
    .Q(\tt_um_rejunity_sn76489.noise[0].gen.lfsr[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17658_ (.D(_00728_),
    .CLK(clknet_leaf_51_clk),
    .Q(\tt_um_rejunity_sn76489.noise[0].gen.lfsr[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17659_ (.D(_00729_),
    .CLK(clknet_leaf_49_clk),
    .Q(\tt_um_rejunity_sn76489.noise[0].gen.lfsr[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17660_ (.D(_00730_),
    .CLK(clknet_leaf_82_clk),
    .Q(\tt_um_rejunity_sn76489.noise[0].gen.counter[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17661_ (.D(_00731_),
    .CLK(clknet_leaf_81_clk),
    .Q(\tt_um_rejunity_sn76489.noise[0].gen.counter[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17662_ (.D(_00732_),
    .CLK(clknet_leaf_58_clk),
    .Q(\tt_um_rejunity_sn76489.noise[0].gen.counter[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17663_ (.D(_00733_),
    .CLK(clknet_leaf_57_clk),
    .Q(\tt_um_rejunity_sn76489.noise[0].gen.counter[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17664_ (.D(_00734_),
    .CLK(clknet_leaf_57_clk),
    .Q(\tt_um_rejunity_sn76489.noise[0].gen.counter[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17665_ (.D(_00735_),
    .CLK(clknet_leaf_57_clk),
    .Q(\tt_um_rejunity_sn76489.noise[0].gen.counter[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17666_ (.D(_00736_),
    .CLK(clknet_leaf_41_clk),
    .Q(\tt_um_rejunity_sn76489.noise[0].gen.counter[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17667_ (.D(_00737_),
    .CLK(clknet_leaf_47_clk),
    .Q(net18));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17668_ (.D(_00738_),
    .CLK(clknet_leaf_80_clk),
    .Q(\tt_um_rejunity_sn76489.tone[2].gen.counter[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17669_ (.D(_00739_),
    .CLK(clknet_leaf_80_clk),
    .Q(\tt_um_rejunity_sn76489.tone[2].gen.counter[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17670_ (.D(_00740_),
    .CLK(clknet_leaf_79_clk),
    .Q(\tt_um_rejunity_sn76489.tone[2].gen.counter[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17671_ (.D(_00741_),
    .CLK(clknet_leaf_79_clk),
    .Q(\tt_um_rejunity_sn76489.tone[2].gen.counter[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17672_ (.D(_00742_),
    .CLK(clknet_leaf_59_clk),
    .Q(\tt_um_rejunity_sn76489.tone[2].gen.counter[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17673_ (.D(_00743_),
    .CLK(clknet_leaf_59_clk),
    .Q(\tt_um_rejunity_sn76489.tone[2].gen.counter[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17674_ (.D(_00744_),
    .CLK(clknet_leaf_81_clk),
    .Q(\tt_um_rejunity_sn76489.tone[2].gen.counter[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17675_ (.D(_00745_),
    .CLK(clknet_leaf_81_clk),
    .Q(\tt_um_rejunity_sn76489.tone[2].gen.counter[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17676_ (.D(_00746_),
    .CLK(clknet_leaf_80_clk),
    .Q(\tt_um_rejunity_sn76489.tone[2].gen.counter[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17677_ (.D(_00747_),
    .CLK(clknet_leaf_61_clk),
    .Q(\tt_um_rejunity_sn76489.tone[2].gen.counter[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17678_ (.D(_00748_),
    .CLK(clknet_leaf_56_clk),
    .Q(\tt_um_rejunity_sn76489.chan[2].attenuation.in ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17679_ (.D(_00749_),
    .CLK(clknet_leaf_68_clk),
    .Q(\tt_um_rejunity_sn76489.tone[1].gen.counter[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17680_ (.D(_00750_),
    .CLK(clknet_leaf_69_clk),
    .Q(\tt_um_rejunity_sn76489.tone[1].gen.counter[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17681_ (.D(_00751_),
    .CLK(clknet_leaf_69_clk),
    .Q(\tt_um_rejunity_sn76489.tone[1].gen.counter[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17682_ (.D(_00752_),
    .CLK(clknet_leaf_70_clk),
    .Q(\tt_um_rejunity_sn76489.tone[1].gen.counter[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17683_ (.D(_00753_),
    .CLK(clknet_leaf_66_clk),
    .Q(\tt_um_rejunity_sn76489.tone[1].gen.counter[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17684_ (.D(_00754_),
    .CLK(clknet_leaf_64_clk),
    .Q(\tt_um_rejunity_sn76489.tone[1].gen.counter[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17685_ (.D(_00755_),
    .CLK(clknet_5_11__leaf_clk),
    .Q(\tt_um_rejunity_sn76489.tone[1].gen.counter[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17686_ (.D(_00756_),
    .CLK(clknet_leaf_66_clk),
    .Q(\tt_um_rejunity_sn76489.tone[1].gen.counter[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17687_ (.D(_00757_),
    .CLK(clknet_leaf_66_clk),
    .Q(\tt_um_rejunity_sn76489.tone[1].gen.counter[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17688_ (.D(_00758_),
    .CLK(clknet_leaf_66_clk),
    .Q(\tt_um_rejunity_sn76489.tone[1].gen.counter[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17689_ (.D(_00759_),
    .CLK(clknet_leaf_63_clk),
    .Q(\tt_um_rejunity_sn76489.chan[1].attenuation.in ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17690_ (.D(_00760_),
    .CLK(clknet_leaf_213_clk),
    .Q(\channels.lfsr[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17691_ (.D(_00761_),
    .CLK(clknet_leaf_216_clk),
    .Q(\channels.lfsr[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17692_ (.D(_00762_),
    .CLK(clknet_leaf_216_clk),
    .Q(\channels.lfsr[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17693_ (.D(_00763_),
    .CLK(clknet_leaf_217_clk),
    .Q(\channels.lfsr[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17694_ (.D(_00764_),
    .CLK(clknet_leaf_220_clk),
    .Q(\channels.lfsr[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17695_ (.D(_00765_),
    .CLK(clknet_leaf_219_clk),
    .Q(\channels.lfsr[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17696_ (.D(_00766_),
    .CLK(clknet_leaf_223_clk),
    .Q(\channels.lfsr[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17697_ (.D(_00767_),
    .CLK(clknet_leaf_221_clk),
    .Q(\channels.lfsr[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17698_ (.D(_00768_),
    .CLK(clknet_leaf_222_clk),
    .Q(\channels.lfsr[0][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17699_ (.D(_00769_),
    .CLK(clknet_leaf_222_clk),
    .Q(\channels.lfsr[0][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17700_ (.D(_00770_),
    .CLK(clknet_leaf_226_clk),
    .Q(\channels.lfsr[0][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17701_ (.D(_00771_),
    .CLK(clknet_leaf_226_clk),
    .Q(\channels.lfsr[0][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17702_ (.D(_00772_),
    .CLK(clknet_leaf_236_clk),
    .Q(\channels.lfsr[0][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17703_ (.D(_00773_),
    .CLK(clknet_leaf_236_clk),
    .Q(\channels.lfsr[0][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17704_ (.D(_00774_),
    .CLK(clknet_leaf_236_clk),
    .Q(\channels.lfsr[0][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17705_ (.D(_00775_),
    .CLK(clknet_leaf_235_clk),
    .Q(\channels.lfsr[0][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17706_ (.D(_00776_),
    .CLK(clknet_leaf_235_clk),
    .Q(\channels.lfsr[0][16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17707_ (.D(_00777_),
    .CLK(clknet_leaf_229_clk),
    .Q(\channels.lfsr[0][17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17708_ (.D(_00778_),
    .CLK(clknet_leaf_229_clk),
    .Q(\channels.lfsr[0][18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17709_ (.D(_00779_),
    .CLK(clknet_leaf_228_clk),
    .Q(\channels.lfsr[0][19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17710_ (.D(_00780_),
    .CLK(clknet_leaf_232_clk),
    .Q(\channels.lfsr[0][20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17711_ (.D(_00781_),
    .CLK(clknet_leaf_231_clk),
    .Q(\channels.lfsr[0][21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17712_ (.D(_00782_),
    .CLK(clknet_leaf_218_clk),
    .Q(\channels.lfsr[0][22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17713_ (.D(_00783_),
    .CLK(clknet_leaf_74_clk),
    .Q(\tt_um_rejunity_sn76489.tone[0].gen.counter[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17714_ (.D(_00784_),
    .CLK(clknet_leaf_67_clk),
    .Q(\tt_um_rejunity_sn76489.tone[0].gen.counter[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17715_ (.D(_00785_),
    .CLK(clknet_leaf_68_clk),
    .Q(\tt_um_rejunity_sn76489.tone[0].gen.counter[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17716_ (.D(_00786_),
    .CLK(clknet_leaf_73_clk),
    .Q(\tt_um_rejunity_sn76489.tone[0].gen.counter[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17717_ (.D(_00787_),
    .CLK(clknet_leaf_67_clk),
    .Q(\tt_um_rejunity_sn76489.tone[0].gen.counter[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17718_ (.D(_00788_),
    .CLK(clknet_leaf_62_clk),
    .Q(\tt_um_rejunity_sn76489.tone[0].gen.counter[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17719_ (.D(_00789_),
    .CLK(clknet_leaf_62_clk),
    .Q(\tt_um_rejunity_sn76489.tone[0].gen.counter[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17720_ (.D(_00790_),
    .CLK(clknet_leaf_67_clk),
    .Q(\tt_um_rejunity_sn76489.tone[0].gen.counter[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17721_ (.D(_00791_),
    .CLK(clknet_leaf_61_clk),
    .Q(\tt_um_rejunity_sn76489.tone[0].gen.counter[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17722_ (.D(_00792_),
    .CLK(clknet_leaf_62_clk),
    .Q(\tt_um_rejunity_sn76489.tone[0].gen.counter[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17723_ (.D(_00793_),
    .CLK(clknet_leaf_53_clk),
    .Q(\tt_um_rejunity_sn76489.chan[0].attenuation.in ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17724_ (.D(_00794_),
    .CLK(clknet_leaf_59_clk),
    .Q(\tt_um_rejunity_sn76489.control_tone_freq[2][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17725_ (.D(_00795_),
    .CLK(clknet_leaf_59_clk),
    .Q(\tt_um_rejunity_sn76489.control_tone_freq[2][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17726_ (.D(_00796_),
    .CLK(clknet_leaf_60_clk),
    .Q(\tt_um_rejunity_sn76489.control_tone_freq[2][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17727_ (.D(_00797_),
    .CLK(clknet_leaf_60_clk),
    .Q(\tt_um_rejunity_sn76489.control_tone_freq[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17728_ (.D(_00798_),
    .CLK(clknet_leaf_60_clk),
    .Q(\tt_um_rejunity_sn76489.control_tone_freq[2][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17729_ (.D(_00799_),
    .CLK(clknet_leaf_60_clk),
    .Q(\tt_um_rejunity_sn76489.control_tone_freq[2][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17730_ (.D(_00800_),
    .CLK(clknet_leaf_64_clk),
    .Q(\tt_um_rejunity_sn76489.control_tone_freq[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17731_ (.D(_00801_),
    .CLK(clknet_leaf_63_clk),
    .Q(\tt_um_rejunity_sn76489.control_tone_freq[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17732_ (.D(_00802_),
    .CLK(clknet_leaf_64_clk),
    .Q(\tt_um_rejunity_sn76489.control_tone_freq[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17733_ (.D(_00803_),
    .CLK(clknet_leaf_64_clk),
    .Q(\tt_um_rejunity_sn76489.control_tone_freq[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17734_ (.D(_00804_),
    .CLK(clknet_leaf_63_clk),
    .Q(\tt_um_rejunity_sn76489.control_tone_freq[1][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17735_ (.D(_00805_),
    .CLK(clknet_leaf_63_clk),
    .Q(\tt_um_rejunity_sn76489.control_tone_freq[1][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17736_ (.D(_00806_),
    .CLK(clknet_leaf_63_clk),
    .Q(\tt_um_rejunity_sn76489.control_tone_freq[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17737_ (.D(_00807_),
    .CLK(clknet_leaf_53_clk),
    .Q(\tt_um_rejunity_sn76489.control_tone_freq[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17738_ (.D(_00808_),
    .CLK(clknet_leaf_53_clk),
    .Q(\tt_um_rejunity_sn76489.control_tone_freq[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17739_ (.D(_00809_),
    .CLK(clknet_leaf_53_clk),
    .Q(\tt_um_rejunity_sn76489.control_tone_freq[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17740_ (.D(_00810_),
    .CLK(clknet_leaf_54_clk),
    .Q(\tt_um_rejunity_sn76489.control_tone_freq[0][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17741_ (.D(_00811_),
    .CLK(clknet_leaf_62_clk),
    .Q(\tt_um_rejunity_sn76489.control_tone_freq[0][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17742_ (.D(_00812_),
    .CLK(clknet_leaf_54_clk),
    .Q(\tt_um_rejunity_sn76489.chan[3].attenuation.control[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17743_ (.D(_00813_),
    .CLK(clknet_leaf_54_clk),
    .Q(\tt_um_rejunity_sn76489.chan[3].attenuation.control[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17744_ (.D(_00814_),
    .CLK(clknet_leaf_54_clk),
    .Q(\tt_um_rejunity_sn76489.chan[3].attenuation.control[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17745_ (.D(_00815_),
    .CLK(clknet_leaf_55_clk),
    .Q(\tt_um_rejunity_sn76489.chan[3].attenuation.control[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17746_ (.D(_00816_),
    .CLK(clknet_leaf_55_clk),
    .Q(\tt_um_rejunity_sn76489.chan[2].attenuation.control[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17747_ (.D(_00817_),
    .CLK(clknet_5_8__leaf_clk),
    .Q(\tt_um_rejunity_sn76489.chan[2].attenuation.control[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17748_ (.D(_00818_),
    .CLK(clknet_leaf_55_clk),
    .Q(\tt_um_rejunity_sn76489.chan[2].attenuation.control[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17749_ (.D(_00819_),
    .CLK(clknet_leaf_55_clk),
    .Q(\tt_um_rejunity_sn76489.chan[2].attenuation.control[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17750_ (.D(_00820_),
    .CLK(clknet_leaf_47_clk),
    .Q(\tt_um_rejunity_sn76489.chan[1].attenuation.control[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17751_ (.D(_00821_),
    .CLK(clknet_leaf_48_clk),
    .Q(\tt_um_rejunity_sn76489.chan[1].attenuation.control[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17752_ (.D(_00822_),
    .CLK(clknet_leaf_48_clk),
    .Q(\tt_um_rejunity_sn76489.chan[1].attenuation.control[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17753_ (.D(_00823_),
    .CLK(clknet_leaf_50_clk),
    .Q(\tt_um_rejunity_sn76489.chan[1].attenuation.control[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17754_ (.D(_00824_),
    .CLK(clknet_leaf_50_clk),
    .Q(\tt_um_rejunity_sn76489.chan[0].attenuation.control[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17755_ (.D(_00825_),
    .CLK(clknet_leaf_49_clk),
    .Q(\tt_um_rejunity_sn76489.chan[0].attenuation.control[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17756_ (.D(_00826_),
    .CLK(clknet_leaf_49_clk),
    .Q(\tt_um_rejunity_sn76489.chan[0].attenuation.control[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17757_ (.D(_00827_),
    .CLK(clknet_leaf_49_clk),
    .Q(\tt_um_rejunity_sn76489.chan[0].attenuation.control[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17758_ (.D(_00828_),
    .CLK(clknet_leaf_81_clk),
    .Q(\tt_um_rejunity_sn76489.noise[0].gen.restart_noise ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17759_ (.D(_00829_),
    .CLK(clknet_leaf_70_clk),
    .Q(\tt_um_rejunity_sn76489.latch_control_reg[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17760_ (.D(_00830_),
    .CLK(clknet_leaf_70_clk),
    .Q(\tt_um_rejunity_sn76489.latch_control_reg[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17761_ (.D(_00831_),
    .CLK(clknet_leaf_70_clk),
    .Q(\tt_um_rejunity_sn76489.latch_control_reg[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17762_ (.D(_00832_),
    .CLK(clknet_5_9__leaf_clk),
    .Q(\tt_um_rejunity_sn76489.clk_counter[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17763_ (.D(_00833_),
    .CLK(clknet_leaf_86_clk),
    .Q(\tt_um_rejunity_sn76489.clk_counter[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17764_ (.D(_00834_),
    .CLK(clknet_leaf_81_clk),
    .Q(\tt_um_rejunity_sn76489.clk_counter[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17765_ (.D(_00835_),
    .CLK(clknet_leaf_82_clk),
    .Q(\tt_um_rejunity_sn76489.clk_counter[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17766_ (.D(_00836_),
    .CLK(clknet_leaf_58_clk),
    .Q(\tt_um_rejunity_sn76489.clk_counter[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17767_ (.D(_00837_),
    .CLK(clknet_leaf_201_clk),
    .Q(\channels.exp_periods[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17768_ (.D(_00838_),
    .CLK(clknet_leaf_203_clk),
    .Q(\channels.exp_periods[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17769_ (.D(_00839_),
    .CLK(clknet_leaf_203_clk),
    .Q(\channels.exp_periods[2][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17770_ (.D(_00840_),
    .CLK(clknet_leaf_201_clk),
    .Q(\channels.exp_periods[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17771_ (.D(_00841_),
    .CLK(clknet_leaf_205_clk),
    .Q(\channels.exp_periods[2][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17772_ (.D(_00842_),
    .CLK(clknet_leaf_200_clk),
    .Q(\channels.exp_periods[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17773_ (.D(_00843_),
    .CLK(clknet_leaf_203_clk),
    .Q(\channels.exp_periods[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17774_ (.D(_00844_),
    .CLK(clknet_leaf_202_clk),
    .Q(\channels.exp_periods[1][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17775_ (.D(_00845_),
    .CLK(clknet_leaf_204_clk),
    .Q(\channels.exp_periods[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17776_ (.D(_00846_),
    .CLK(clknet_leaf_206_clk),
    .Q(\channels.exp_periods[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17777_ (.D(_00847_),
    .CLK(clknet_leaf_195_clk),
    .Q(\channels.exp_counter[3][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17778_ (.D(_00848_),
    .CLK(clknet_leaf_196_clk),
    .Q(\channels.exp_counter[3][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17779_ (.D(_00849_),
    .CLK(clknet_leaf_197_clk),
    .Q(\channels.exp_counter[3][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17780_ (.D(_00850_),
    .CLK(clknet_leaf_197_clk),
    .Q(\channels.exp_counter[3][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17781_ (.D(_00851_),
    .CLK(clknet_leaf_206_clk),
    .Q(\channels.exp_counter[3][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17782_ (.D(_00852_),
    .CLK(clknet_leaf_200_clk),
    .Q(\channels.exp_periods[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17783_ (.D(_00853_),
    .CLK(clknet_leaf_214_clk),
    .Q(\channels.exp_periods[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17784_ (.D(_00854_),
    .CLK(clknet_leaf_215_clk),
    .Q(\channels.exp_periods[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17785_ (.D(_00855_),
    .CLK(clknet_leaf_204_clk),
    .Q(\channels.exp_periods[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17786_ (.D(_00856_),
    .CLK(clknet_leaf_205_clk),
    .Q(\channels.exp_periods[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17787_ (.D(_00857_),
    .CLK(clknet_leaf_56_clk),
    .Q(\tt_um_rejunity_sn76489.control_noise[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17788_ (.D(_00858_),
    .CLK(clknet_leaf_56_clk),
    .Q(\tt_um_rejunity_sn76489.control_noise[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17789_ (.D(_00859_),
    .CLK(clknet_leaf_49_clk),
    .Q(\tt_um_rejunity_sn76489.control_noise[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_0_clk (.I(clk),
    .Z(clknet_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_0_0_clk (.I(clknet_0_clk),
    .Z(clknet_3_0_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_1_0_clk (.I(clknet_0_clk),
    .Z(clknet_3_1_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_2_0_clk (.I(clknet_0_clk),
    .Z(clknet_3_2_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_3_0_clk (.I(clknet_0_clk),
    .Z(clknet_3_3_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_4_0_clk (.I(clknet_0_clk),
    .Z(clknet_3_4_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_5_0_clk (.I(clknet_0_clk),
    .Z(clknet_3_5_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_6_0_clk (.I(clknet_0_clk),
    .Z(clknet_3_6_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_7_0_clk (.I(clknet_0_clk),
    .Z(clknet_3_7_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_5_0__f_clk (.I(clknet_3_0_0_clk),
    .Z(clknet_5_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_5_10__f_clk (.I(clknet_3_2_0_clk),
    .Z(clknet_5_10__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_5_11__f_clk (.I(clknet_3_2_0_clk),
    .Z(clknet_5_11__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_5_12__f_clk (.I(clknet_3_3_0_clk),
    .Z(clknet_5_12__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_5_13__f_clk (.I(clknet_3_3_0_clk),
    .Z(clknet_5_13__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_5_14__f_clk (.I(clknet_3_3_0_clk),
    .Z(clknet_5_14__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_5_15__f_clk (.I(clknet_3_3_0_clk),
    .Z(clknet_5_15__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_5_16__f_clk (.I(clknet_3_4_0_clk),
    .Z(clknet_5_16__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_5_17__f_clk (.I(clknet_3_4_0_clk),
    .Z(clknet_5_17__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_5_18__f_clk (.I(clknet_3_4_0_clk),
    .Z(clknet_5_18__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_5_19__f_clk (.I(clknet_3_4_0_clk),
    .Z(clknet_5_19__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_5_1__f_clk (.I(clknet_3_0_0_clk),
    .Z(clknet_5_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_5_20__f_clk (.I(clknet_3_5_0_clk),
    .Z(clknet_5_20__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_5_21__f_clk (.I(clknet_3_5_0_clk),
    .Z(clknet_5_21__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_5_22__f_clk (.I(clknet_3_5_0_clk),
    .Z(clknet_5_22__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_5_23__f_clk (.I(clknet_3_5_0_clk),
    .Z(clknet_5_23__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_5_24__f_clk (.I(clknet_3_6_0_clk),
    .Z(clknet_5_24__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_5_25__f_clk (.I(clknet_3_6_0_clk),
    .Z(clknet_5_25__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_5_26__f_clk (.I(clknet_3_6_0_clk),
    .Z(clknet_5_26__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_5_27__f_clk (.I(clknet_3_6_0_clk),
    .Z(clknet_5_27__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_5_28__f_clk (.I(clknet_3_7_0_clk),
    .Z(clknet_5_28__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_5_29__f_clk (.I(clknet_3_7_0_clk),
    .Z(clknet_5_29__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_5_2__f_clk (.I(clknet_3_0_0_clk),
    .Z(clknet_5_2__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_5_30__f_clk (.I(clknet_3_7_0_clk),
    .Z(clknet_5_30__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_5_31__f_clk (.I(clknet_3_7_0_clk),
    .Z(clknet_5_31__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_5_3__f_clk (.I(clknet_3_0_0_clk),
    .Z(clknet_5_3__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_5_4__f_clk (.I(clknet_3_1_0_clk),
    .Z(clknet_5_4__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_5_5__f_clk (.I(clknet_3_1_0_clk),
    .Z(clknet_5_5__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_5_6__f_clk (.I(clknet_3_1_0_clk),
    .Z(clknet_5_6__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_5_7__f_clk (.I(clknet_3_1_0_clk),
    .Z(clknet_5_7__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_5_8__f_clk (.I(clknet_3_2_0_clk),
    .Z(clknet_5_8__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_5_9__f_clk (.I(clknet_3_2_0_clk),
    .Z(clknet_5_9__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_0_clk (.I(clknet_5_4__leaf_clk),
    .Z(clknet_leaf_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_100_clk (.I(clknet_5_13__leaf_clk),
    .Z(clknet_leaf_100_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_101_clk (.I(clknet_5_13__leaf_clk),
    .Z(clknet_leaf_101_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_102_clk (.I(clknet_5_13__leaf_clk),
    .Z(clknet_leaf_102_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_103_clk (.I(clknet_5_13__leaf_clk),
    .Z(clknet_leaf_103_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_104_clk (.I(clknet_5_13__leaf_clk),
    .Z(clknet_leaf_104_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_105_clk (.I(clknet_5_15__leaf_clk),
    .Z(clknet_leaf_105_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_106_clk (.I(clknet_5_15__leaf_clk),
    .Z(clknet_leaf_106_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_107_clk (.I(clknet_5_15__leaf_clk),
    .Z(clknet_leaf_107_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_108_clk (.I(clknet_5_15__leaf_clk),
    .Z(clknet_leaf_108_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_109_clk (.I(clknet_5_15__leaf_clk),
    .Z(clknet_leaf_109_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_110_clk (.I(clknet_5_15__leaf_clk),
    .Z(clknet_leaf_110_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_111_clk (.I(clknet_5_15__leaf_clk),
    .Z(clknet_leaf_111_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_112_clk (.I(clknet_5_15__leaf_clk),
    .Z(clknet_leaf_112_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_113_clk (.I(clknet_5_15__leaf_clk),
    .Z(clknet_leaf_113_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_114_clk (.I(clknet_5_26__leaf_clk),
    .Z(clknet_leaf_114_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_115_clk (.I(clknet_5_26__leaf_clk),
    .Z(clknet_leaf_115_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_116_clk (.I(clknet_5_26__leaf_clk),
    .Z(clknet_leaf_116_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_117_clk (.I(clknet_5_27__leaf_clk),
    .Z(clknet_leaf_117_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_118_clk (.I(clknet_5_26__leaf_clk),
    .Z(clknet_leaf_118_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_119_clk (.I(clknet_5_26__leaf_clk),
    .Z(clknet_leaf_119_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_11_clk (.I(clknet_5_7__leaf_clk),
    .Z(clknet_leaf_11_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_121_clk (.I(clknet_5_27__leaf_clk),
    .Z(clknet_leaf_121_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_122_clk (.I(clknet_5_30__leaf_clk),
    .Z(clknet_leaf_122_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_123_clk (.I(clknet_5_30__leaf_clk),
    .Z(clknet_leaf_123_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_124_clk (.I(clknet_5_27__leaf_clk),
    .Z(clknet_leaf_124_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_125_clk (.I(clknet_5_27__leaf_clk),
    .Z(clknet_leaf_125_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_127_clk (.I(clknet_5_27__leaf_clk),
    .Z(clknet_leaf_127_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_128_clk (.I(clknet_5_30__leaf_clk),
    .Z(clknet_leaf_128_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_129_clk (.I(clknet_5_30__leaf_clk),
    .Z(clknet_leaf_129_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_130_clk (.I(clknet_5_30__leaf_clk),
    .Z(clknet_leaf_130_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_131_clk (.I(clknet_5_31__leaf_clk),
    .Z(clknet_leaf_131_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_132_clk (.I(clknet_5_31__leaf_clk),
    .Z(clknet_leaf_132_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_133_clk (.I(clknet_5_31__leaf_clk),
    .Z(clknet_leaf_133_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_134_clk (.I(clknet_5_31__leaf_clk),
    .Z(clknet_leaf_134_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_135_clk (.I(clknet_5_31__leaf_clk),
    .Z(clknet_leaf_135_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_136_clk (.I(clknet_5_31__leaf_clk),
    .Z(clknet_leaf_136_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_137_clk (.I(clknet_5_31__leaf_clk),
    .Z(clknet_leaf_137_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_138_clk (.I(clknet_5_31__leaf_clk),
    .Z(clknet_leaf_138_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_139_clk (.I(clknet_5_31__leaf_clk),
    .Z(clknet_leaf_139_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_13_clk (.I(clknet_5_6__leaf_clk),
    .Z(clknet_leaf_13_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_141_clk (.I(clknet_5_30__leaf_clk),
    .Z(clknet_leaf_141_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_142_clk (.I(clknet_5_30__leaf_clk),
    .Z(clknet_leaf_142_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_143_clk (.I(clknet_5_27__leaf_clk),
    .Z(clknet_leaf_143_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_144_clk (.I(clknet_5_30__leaf_clk),
    .Z(clknet_leaf_144_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_145_clk (.I(clknet_5_30__leaf_clk),
    .Z(clknet_leaf_145_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_146_clk (.I(clknet_5_28__leaf_clk),
    .Z(clknet_leaf_146_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_147_clk (.I(clknet_5_29__leaf_clk),
    .Z(clknet_leaf_147_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_148_clk (.I(clknet_5_31__leaf_clk),
    .Z(clknet_leaf_148_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_149_clk (.I(clknet_5_31__leaf_clk),
    .Z(clknet_leaf_149_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_14_clk (.I(clknet_5_6__leaf_clk),
    .Z(clknet_leaf_14_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_150_clk (.I(clknet_5_29__leaf_clk),
    .Z(clknet_leaf_150_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_151_clk (.I(clknet_5_29__leaf_clk),
    .Z(clknet_leaf_151_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_152_clk (.I(clknet_5_29__leaf_clk),
    .Z(clknet_leaf_152_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_153_clk (.I(clknet_5_29__leaf_clk),
    .Z(clknet_leaf_153_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_154_clk (.I(clknet_5_29__leaf_clk),
    .Z(clknet_leaf_154_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_155_clk (.I(clknet_5_29__leaf_clk),
    .Z(clknet_leaf_155_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_156_clk (.I(clknet_5_29__leaf_clk),
    .Z(clknet_leaf_156_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_157_clk (.I(clknet_5_29__leaf_clk),
    .Z(clknet_leaf_157_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_158_clk (.I(clknet_5_28__leaf_clk),
    .Z(clknet_leaf_158_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_159_clk (.I(clknet_5_28__leaf_clk),
    .Z(clknet_leaf_159_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_15_clk (.I(clknet_5_6__leaf_clk),
    .Z(clknet_leaf_15_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_161_clk (.I(clknet_5_28__leaf_clk),
    .Z(clknet_leaf_161_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_162_clk (.I(clknet_5_25__leaf_clk),
    .Z(clknet_leaf_162_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_163_clk (.I(clknet_5_28__leaf_clk),
    .Z(clknet_leaf_163_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_164_clk (.I(clknet_5_28__leaf_clk),
    .Z(clknet_leaf_164_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_165_clk (.I(clknet_5_25__leaf_clk),
    .Z(clknet_leaf_165_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_166_clk (.I(clknet_5_25__leaf_clk),
    .Z(clknet_leaf_166_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_168_clk (.I(clknet_5_25__leaf_clk),
    .Z(clknet_leaf_168_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_169_clk (.I(clknet_5_24__leaf_clk),
    .Z(clknet_leaf_169_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_170_clk (.I(clknet_5_24__leaf_clk),
    .Z(clknet_leaf_170_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_171_clk (.I(clknet_5_24__leaf_clk),
    .Z(clknet_leaf_171_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_172_clk (.I(clknet_5_24__leaf_clk),
    .Z(clknet_leaf_172_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_173_clk (.I(clknet_5_24__leaf_clk),
    .Z(clknet_leaf_173_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_174_clk (.I(clknet_5_24__leaf_clk),
    .Z(clknet_leaf_174_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_175_clk (.I(clknet_5_18__leaf_clk),
    .Z(clknet_leaf_175_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_176_clk (.I(clknet_5_18__leaf_clk),
    .Z(clknet_leaf_176_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_177_clk (.I(clknet_5_18__leaf_clk),
    .Z(clknet_leaf_177_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_178_clk (.I(clknet_5_18__leaf_clk),
    .Z(clknet_leaf_178_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_179_clk (.I(clknet_5_18__leaf_clk),
    .Z(clknet_leaf_179_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_180_clk (.I(clknet_5_19__leaf_clk),
    .Z(clknet_leaf_180_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_181_clk (.I(clknet_5_19__leaf_clk),
    .Z(clknet_leaf_181_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_182_clk (.I(clknet_5_19__leaf_clk),
    .Z(clknet_leaf_182_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_185_clk (.I(clknet_5_22__leaf_clk),
    .Z(clknet_leaf_185_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_186_clk (.I(clknet_5_22__leaf_clk),
    .Z(clknet_leaf_186_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_187_clk (.I(clknet_5_19__leaf_clk),
    .Z(clknet_leaf_187_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_188_clk (.I(clknet_5_19__leaf_clk),
    .Z(clknet_leaf_188_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_189_clk (.I(clknet_5_22__leaf_clk),
    .Z(clknet_leaf_189_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_18_clk (.I(clknet_5_6__leaf_clk),
    .Z(clknet_leaf_18_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_190_clk (.I(clknet_5_22__leaf_clk),
    .Z(clknet_leaf_190_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_191_clk (.I(clknet_5_22__leaf_clk),
    .Z(clknet_leaf_191_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_192_clk (.I(clknet_5_23__leaf_clk),
    .Z(clknet_leaf_192_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_193_clk (.I(clknet_5_23__leaf_clk),
    .Z(clknet_leaf_193_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_194_clk (.I(clknet_5_23__leaf_clk),
    .Z(clknet_leaf_194_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_195_clk (.I(clknet_5_23__leaf_clk),
    .Z(clknet_leaf_195_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_196_clk (.I(clknet_5_23__leaf_clk),
    .Z(clknet_leaf_196_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_197_clk (.I(clknet_5_23__leaf_clk),
    .Z(clknet_leaf_197_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_19_clk (.I(clknet_5_3__leaf_clk),
    .Z(clknet_leaf_19_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_1_clk (.I(clknet_5_4__leaf_clk),
    .Z(clknet_leaf_1_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_200_clk (.I(clknet_5_23__leaf_clk),
    .Z(clknet_leaf_200_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_201_clk (.I(clknet_5_23__leaf_clk),
    .Z(clknet_leaf_201_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_202_clk (.I(clknet_5_21__leaf_clk),
    .Z(clknet_leaf_202_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_203_clk (.I(clknet_5_21__leaf_clk),
    .Z(clknet_leaf_203_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_204_clk (.I(clknet_5_22__leaf_clk),
    .Z(clknet_leaf_204_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_205_clk (.I(clknet_5_23__leaf_clk),
    .Z(clknet_leaf_205_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_206_clk (.I(clknet_5_22__leaf_clk),
    .Z(clknet_leaf_206_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_207_clk (.I(clknet_5_20__leaf_clk),
    .Z(clknet_leaf_207_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_208_clk (.I(clknet_5_22__leaf_clk),
    .Z(clknet_leaf_208_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_209_clk (.I(clknet_5_17__leaf_clk),
    .Z(clknet_leaf_209_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_20_clk (.I(clknet_5_3__leaf_clk),
    .Z(clknet_leaf_20_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_210_clk (.I(clknet_5_20__leaf_clk),
    .Z(clknet_leaf_210_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_211_clk (.I(clknet_5_20__leaf_clk),
    .Z(clknet_leaf_211_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_212_clk (.I(clknet_5_20__leaf_clk),
    .Z(clknet_leaf_212_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_213_clk (.I(clknet_5_21__leaf_clk),
    .Z(clknet_leaf_213_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_214_clk (.I(clknet_5_21__leaf_clk),
    .Z(clknet_leaf_214_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_215_clk (.I(clknet_5_21__leaf_clk),
    .Z(clknet_leaf_215_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_216_clk (.I(clknet_5_21__leaf_clk),
    .Z(clknet_leaf_216_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_217_clk (.I(clknet_5_21__leaf_clk),
    .Z(clknet_leaf_217_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_218_clk (.I(clknet_5_21__leaf_clk),
    .Z(clknet_leaf_218_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_219_clk (.I(clknet_5_21__leaf_clk),
    .Z(clknet_leaf_219_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_21_clk (.I(clknet_5_3__leaf_clk),
    .Z(clknet_leaf_21_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_220_clk (.I(clknet_5_21__leaf_clk),
    .Z(clknet_leaf_220_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_221_clk (.I(clknet_5_21__leaf_clk),
    .Z(clknet_leaf_221_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_222_clk (.I(clknet_5_20__leaf_clk),
    .Z(clknet_leaf_222_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_223_clk (.I(clknet_5_20__leaf_clk),
    .Z(clknet_leaf_223_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_224_clk (.I(clknet_5_20__leaf_clk),
    .Z(clknet_leaf_224_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_225_clk (.I(clknet_5_20__leaf_clk),
    .Z(clknet_leaf_225_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_226_clk (.I(clknet_5_20__leaf_clk),
    .Z(clknet_leaf_226_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_227_clk (.I(clknet_5_17__leaf_clk),
    .Z(clknet_leaf_227_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_228_clk (.I(clknet_5_17__leaf_clk),
    .Z(clknet_leaf_228_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_229_clk (.I(clknet_5_17__leaf_clk),
    .Z(clknet_leaf_229_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_22_clk (.I(clknet_5_3__leaf_clk),
    .Z(clknet_leaf_22_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_230_clk (.I(clknet_5_17__leaf_clk),
    .Z(clknet_leaf_230_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_231_clk (.I(clknet_5_20__leaf_clk),
    .Z(clknet_leaf_231_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_232_clk (.I(clknet_5_17__leaf_clk),
    .Z(clknet_leaf_232_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_233_clk (.I(clknet_5_17__leaf_clk),
    .Z(clknet_leaf_233_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_235_clk (.I(clknet_5_16__leaf_clk),
    .Z(clknet_leaf_235_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_236_clk (.I(clknet_5_16__leaf_clk),
    .Z(clknet_leaf_236_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_238_clk (.I(clknet_5_16__leaf_clk),
    .Z(clknet_leaf_238_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_239_clk (.I(clknet_5_16__leaf_clk),
    .Z(clknet_leaf_239_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_23_clk (.I(clknet_5_1__leaf_clk),
    .Z(clknet_leaf_23_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_240_clk (.I(clknet_5_18__leaf_clk),
    .Z(clknet_leaf_240_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_242_clk (.I(clknet_5_18__leaf_clk),
    .Z(clknet_leaf_242_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_243_clk (.I(clknet_5_5__leaf_clk),
    .Z(clknet_leaf_243_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_244_clk (.I(clknet_5_0__leaf_clk),
    .Z(clknet_leaf_244_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_245_clk (.I(clknet_5_0__leaf_clk),
    .Z(clknet_leaf_245_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_246_clk (.I(clknet_5_0__leaf_clk),
    .Z(clknet_leaf_246_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_247_clk (.I(clknet_5_0__leaf_clk),
    .Z(clknet_leaf_247_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_248_clk (.I(clknet_5_1__leaf_clk),
    .Z(clknet_leaf_248_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_249_clk (.I(clknet_5_1__leaf_clk),
    .Z(clknet_leaf_249_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_25_clk (.I(clknet_5_6__leaf_clk),
    .Z(clknet_leaf_25_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_26_clk (.I(clknet_5_4__leaf_clk),
    .Z(clknet_leaf_26_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_27_clk (.I(clknet_5_1__leaf_clk),
    .Z(clknet_leaf_27_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_29_clk (.I(clknet_5_0__leaf_clk),
    .Z(clknet_leaf_29_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_2_clk (.I(clknet_5_1__leaf_clk),
    .Z(clknet_leaf_2_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_30_clk (.I(clknet_5_0__leaf_clk),
    .Z(clknet_leaf_30_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_32_clk (.I(clknet_5_2__leaf_clk),
    .Z(clknet_leaf_32_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_33_clk (.I(clknet_5_2__leaf_clk),
    .Z(clknet_leaf_33_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_34_clk (.I(clknet_5_2__leaf_clk),
    .Z(clknet_leaf_34_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_37_clk (.I(clknet_5_3__leaf_clk),
    .Z(clknet_leaf_37_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_38_clk (.I(clknet_5_3__leaf_clk),
    .Z(clknet_leaf_38_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_39_clk (.I(clknet_5_3__leaf_clk),
    .Z(clknet_leaf_39_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_40_clk (.I(clknet_5_3__leaf_clk),
    .Z(clknet_leaf_40_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_41_clk (.I(clknet_5_3__leaf_clk),
    .Z(clknet_leaf_41_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_42_clk (.I(clknet_5_3__leaf_clk),
    .Z(clknet_leaf_42_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_44_clk (.I(clknet_5_2__leaf_clk),
    .Z(clknet_leaf_44_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_45_clk (.I(clknet_5_2__leaf_clk),
    .Z(clknet_leaf_45_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_46_clk (.I(clknet_5_2__leaf_clk),
    .Z(clknet_leaf_46_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_47_clk (.I(clknet_5_10__leaf_clk),
    .Z(clknet_leaf_47_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_48_clk (.I(clknet_5_10__leaf_clk),
    .Z(clknet_leaf_48_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_49_clk (.I(clknet_5_10__leaf_clk),
    .Z(clknet_leaf_49_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_4_clk (.I(clknet_5_4__leaf_clk),
    .Z(clknet_leaf_4_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_50_clk (.I(clknet_5_10__leaf_clk),
    .Z(clknet_leaf_50_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_51_clk (.I(clknet_5_10__leaf_clk),
    .Z(clknet_leaf_51_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_52_clk (.I(clknet_5_10__leaf_clk),
    .Z(clknet_leaf_52_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_53_clk (.I(clknet_5_10__leaf_clk),
    .Z(clknet_leaf_53_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_54_clk (.I(clknet_5_10__leaf_clk),
    .Z(clknet_leaf_54_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_55_clk (.I(clknet_5_8__leaf_clk),
    .Z(clknet_leaf_55_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_56_clk (.I(clknet_5_8__leaf_clk),
    .Z(clknet_leaf_56_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_57_clk (.I(clknet_5_3__leaf_clk),
    .Z(clknet_leaf_57_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_58_clk (.I(clknet_5_8__leaf_clk),
    .Z(clknet_leaf_58_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_59_clk (.I(clknet_5_8__leaf_clk),
    .Z(clknet_leaf_59_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_5_clk (.I(clknet_5_4__leaf_clk),
    .Z(clknet_leaf_5_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_60_clk (.I(clknet_5_8__leaf_clk),
    .Z(clknet_leaf_60_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_61_clk (.I(clknet_5_9__leaf_clk),
    .Z(clknet_leaf_61_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_62_clk (.I(clknet_5_11__leaf_clk),
    .Z(clknet_leaf_62_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_63_clk (.I(clknet_5_11__leaf_clk),
    .Z(clknet_leaf_63_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_64_clk (.I(clknet_5_11__leaf_clk),
    .Z(clknet_leaf_64_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_66_clk (.I(clknet_5_11__leaf_clk),
    .Z(clknet_leaf_66_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_67_clk (.I(clknet_5_11__leaf_clk),
    .Z(clknet_leaf_67_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_68_clk (.I(clknet_5_11__leaf_clk),
    .Z(clknet_leaf_68_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_69_clk (.I(clknet_5_11__leaf_clk),
    .Z(clknet_leaf_69_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_6_clk (.I(clknet_5_5__leaf_clk),
    .Z(clknet_leaf_6_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_70_clk (.I(clknet_5_14__leaf_clk),
    .Z(clknet_leaf_70_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_71_clk (.I(clknet_5_14__leaf_clk),
    .Z(clknet_leaf_71_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_72_clk (.I(clknet_5_14__leaf_clk),
    .Z(clknet_leaf_72_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_73_clk (.I(clknet_5_14__leaf_clk),
    .Z(clknet_leaf_73_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_74_clk (.I(clknet_5_9__leaf_clk),
    .Z(clknet_leaf_74_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_75_clk (.I(clknet_5_14__leaf_clk),
    .Z(clknet_leaf_75_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_76_clk (.I(clknet_5_14__leaf_clk),
    .Z(clknet_leaf_76_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_77_clk (.I(clknet_5_12__leaf_clk),
    .Z(clknet_leaf_77_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_78_clk (.I(clknet_5_12__leaf_clk),
    .Z(clknet_leaf_78_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_79_clk (.I(clknet_5_12__leaf_clk),
    .Z(clknet_leaf_79_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_80_clk (.I(clknet_5_9__leaf_clk),
    .Z(clknet_leaf_80_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_81_clk (.I(clknet_5_9__leaf_clk),
    .Z(clknet_leaf_81_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_82_clk (.I(clknet_5_9__leaf_clk),
    .Z(clknet_leaf_82_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_85_clk (.I(clknet_5_12__leaf_clk),
    .Z(clknet_leaf_85_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_86_clk (.I(clknet_5_12__leaf_clk),
    .Z(clknet_leaf_86_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_87_clk (.I(clknet_5_12__leaf_clk),
    .Z(clknet_leaf_87_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_88_clk (.I(clknet_5_12__leaf_clk),
    .Z(clknet_leaf_88_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_89_clk (.I(clknet_5_12__leaf_clk),
    .Z(clknet_leaf_89_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_8_clk (.I(clknet_5_5__leaf_clk),
    .Z(clknet_leaf_8_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_90_clk (.I(clknet_5_12__leaf_clk),
    .Z(clknet_leaf_90_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_91_clk (.I(clknet_5_7__leaf_clk),
    .Z(clknet_leaf_91_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_93_clk (.I(clknet_5_7__leaf_clk),
    .Z(clknet_leaf_93_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_94_clk (.I(clknet_5_7__leaf_clk),
    .Z(clknet_leaf_94_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_95_clk (.I(clknet_5_13__leaf_clk),
    .Z(clknet_leaf_95_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_96_clk (.I(clknet_5_13__leaf_clk),
    .Z(clknet_leaf_96_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_97_clk (.I(clknet_5_13__leaf_clk),
    .Z(clknet_leaf_97_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_98_clk (.I(clknet_5_13__leaf_clk),
    .Z(clknet_leaf_98_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_99_clk (.I(clknet_5_13__leaf_clk),
    .Z(clknet_leaf_99_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_9_clk (.I(clknet_5_5__leaf_clk),
    .Z(clknet_leaf_9_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 input1 (.I(addr[0]),
    .Z(net1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input10 (.I(bus_in[2]),
    .Z(net10));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input11 (.I(bus_in[3]),
    .Z(net11));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input12 (.I(bus_in[4]),
    .Z(net12));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input13 (.I(bus_in[5]),
    .Z(net13));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input14 (.I(bus_in[6]),
    .Z(net14));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input15 (.I(bus_in[7]),
    .Z(net15));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input16 (.I(bus_we),
    .Z(net16));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 input17 (.I(rst),
    .Z(net17));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input2 (.I(addr[1]),
    .Z(net2));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 input3 (.I(addr[2]),
    .Z(net3));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input4 (.I(addr[3]),
    .Z(net4));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input5 (.I(addr[4]),
    .Z(net5));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input6 (.I(addr[5]),
    .Z(net6));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input7 (.I(bus_cyc),
    .Z(net7));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input8 (.I(bus_in[0]),
    .Z(net8));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input9 (.I(bus_in[1]),
    .Z(net9));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output18 (.I(net18),
    .Z(DAC_clk));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output19 (.I(net19),
    .Z(DAC_dat_1));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output20 (.I(net20),
    .Z(DAC_dat_2));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output21 (.I(net21),
    .Z(DAC_le));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output22 (.I(net22),
    .Z(bus_out[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output23 (.I(net23),
    .Z(bus_out[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output24 (.I(net24),
    .Z(bus_out[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output25 (.I(net25),
    .Z(bus_out[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output26 (.I(net26),
    .Z(bus_out[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output27 (.I(net27),
    .Z(bus_out[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output28 (.I(net28),
    .Z(bus_out[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output29 (.I(net29),
    .Z(bus_out[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 rebuffer1 (.I(net43),
    .Z(net30));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer10 (.I(_05431_),
    .Z(net39));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer11 (.I(_05431_),
    .Z(net40));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer12 (.I(_05060_),
    .Z(net41));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer13 (.I(net53),
    .Z(net42));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer14 (.I(_06709_),
    .Z(net43));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer15 (.I(_05375_),
    .Z(net44));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 rebuffer16 (.I(_05287_),
    .Z(net45));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 rebuffer17 (.I(_06063_),
    .Z(net46));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer18 (.I(_05330_),
    .Z(net47));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer19 (.I(_05182_),
    .Z(net48));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 rebuffer2 (.I(_05037_),
    .Z(net31));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer20 (.I(_05151_),
    .Z(net49));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer21 (.I(_04812_),
    .Z(net50));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer22 (.I(_06304_),
    .Z(net51));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer23 (.I(_04988_),
    .Z(net52));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer24 (.I(net54),
    .Z(net53));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 rebuffer25 (.I(net65),
    .Z(net54));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 rebuffer26 (.I(_05378_),
    .Z(net55));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer27 (.I(net55),
    .Z(net56));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer28 (.I(_04235_),
    .Z(net57));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer29 (.I(_04880_),
    .Z(net58));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 rebuffer3 (.I(net42),
    .Z(net32));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer30 (.I(_04162_),
    .Z(net59));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 rebuffer31 (.I(_04177_),
    .Z(net60));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer32 (.I(_05411_),
    .Z(net61));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer33 (.I(_05475_),
    .Z(net62));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer34 (.I(_03286_),
    .Z(net63));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer35 (.I(net63),
    .Z(net64));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 rebuffer36 (.I(_06835_),
    .Z(net65));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 rebuffer37 (.I(_05413_),
    .Z(net66));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer38 (.I(_07426_),
    .Z(net67));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer39 (.I(_04388_),
    .Z(net68));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer4 (.I(_04409_),
    .Z(net33));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer40 (.I(_05228_),
    .Z(net69));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer41 (.I(_06896_),
    .Z(net70));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 rebuffer42 (.I(_04493_),
    .Z(net71));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer5 (.I(_04346_),
    .Z(net34));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 rebuffer6 (.I(_05423_),
    .Z(net35));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer7 (.I(_07362_),
    .Z(net36));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer8 (.I(_05031_),
    .Z(net37));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer9 (.I(net37),
    .Z(net38));
endmodule

