magic
tech gf180mcuC
magscale 1 5
timestamp 1684423258
<< obsm1 >>
rect 118172 170471 206820 227561
<< metal2 >>
rect 5516 297780 5628 298500
rect 16548 297780 16660 298500
rect 27580 297780 27692 298500
rect 38612 297780 38724 298500
rect 49644 297780 49756 298500
rect 60676 297780 60788 298500
rect 71708 297780 71820 298500
rect 82740 297780 82852 298500
rect 93772 297780 93884 298500
rect 104804 297780 104916 298500
rect 115836 297780 115948 298500
rect 126868 297780 126980 298500
rect 137900 297780 138012 298500
rect 148932 297780 149044 298500
rect 159964 297780 160076 298500
rect 170996 297780 171108 298500
rect 182028 297780 182140 298500
rect 193060 297780 193172 298500
rect 204092 297780 204204 298500
rect 215124 297780 215236 298500
rect 226156 297780 226268 298500
rect 237188 297780 237300 298500
rect 248220 297780 248332 298500
rect 259252 297780 259364 298500
rect 270284 297780 270396 298500
rect 281316 297780 281428 298500
rect 292348 297780 292460 298500
rect 5684 -480 5796 240
rect 6636 -480 6748 240
rect 7588 -480 7700 240
rect 8540 -480 8652 240
rect 9492 -480 9604 240
rect 10444 -480 10556 240
rect 11396 -480 11508 240
rect 12348 -480 12460 240
rect 13300 -480 13412 240
rect 14252 -480 14364 240
rect 15204 -480 15316 240
rect 16156 -480 16268 240
rect 17108 -480 17220 240
rect 18060 -480 18172 240
rect 19012 -480 19124 240
rect 19964 -480 20076 240
rect 20916 -480 21028 240
rect 21868 -480 21980 240
rect 22820 -480 22932 240
rect 23772 -480 23884 240
rect 24724 -480 24836 240
rect 25676 -480 25788 240
rect 26628 -480 26740 240
rect 27580 -480 27692 240
rect 28532 -480 28644 240
rect 29484 -480 29596 240
rect 30436 -480 30548 240
rect 31388 -480 31500 240
rect 32340 -480 32452 240
rect 33292 -480 33404 240
rect 34244 -480 34356 240
rect 35196 -480 35308 240
rect 36148 -480 36260 240
rect 37100 -480 37212 240
rect 38052 -480 38164 240
rect 39004 -480 39116 240
rect 39956 -480 40068 240
rect 40908 -480 41020 240
rect 41860 -480 41972 240
rect 42812 -480 42924 240
rect 43764 -480 43876 240
rect 44716 -480 44828 240
rect 45668 -480 45780 240
rect 46620 -480 46732 240
rect 47572 -480 47684 240
rect 48524 -480 48636 240
rect 49476 -480 49588 240
rect 50428 -480 50540 240
rect 51380 -480 51492 240
rect 52332 -480 52444 240
rect 53284 -480 53396 240
rect 54236 -480 54348 240
rect 55188 -480 55300 240
rect 56140 -480 56252 240
rect 57092 -480 57204 240
rect 58044 -480 58156 240
rect 58996 -480 59108 240
rect 59948 -480 60060 240
rect 60900 -480 61012 240
rect 61852 -480 61964 240
rect 62804 -480 62916 240
rect 63756 -480 63868 240
rect 64708 -480 64820 240
rect 65660 -480 65772 240
rect 66612 -480 66724 240
rect 67564 -480 67676 240
rect 68516 -480 68628 240
rect 69468 -480 69580 240
rect 70420 -480 70532 240
rect 71372 -480 71484 240
rect 72324 -480 72436 240
rect 73276 -480 73388 240
rect 74228 -480 74340 240
rect 75180 -480 75292 240
rect 76132 -480 76244 240
rect 77084 -480 77196 240
rect 78036 -480 78148 240
rect 78988 -480 79100 240
rect 79940 -480 80052 240
rect 80892 -480 81004 240
rect 81844 -480 81956 240
rect 82796 -480 82908 240
rect 83748 -480 83860 240
rect 84700 -480 84812 240
rect 85652 -480 85764 240
rect 86604 -480 86716 240
rect 87556 -480 87668 240
rect 88508 -480 88620 240
rect 89460 -480 89572 240
rect 90412 -480 90524 240
rect 91364 -480 91476 240
rect 92316 -480 92428 240
rect 93268 -480 93380 240
rect 94220 -480 94332 240
rect 95172 -480 95284 240
rect 96124 -480 96236 240
rect 97076 -480 97188 240
rect 98028 -480 98140 240
rect 98980 -480 99092 240
rect 99932 -480 100044 240
rect 100884 -480 100996 240
rect 101836 -480 101948 240
rect 102788 -480 102900 240
rect 103740 -480 103852 240
rect 104692 -480 104804 240
rect 105644 -480 105756 240
rect 106596 -480 106708 240
rect 107548 -480 107660 240
rect 108500 -480 108612 240
rect 109452 -480 109564 240
rect 110404 -480 110516 240
rect 111356 -480 111468 240
rect 112308 -480 112420 240
rect 113260 -480 113372 240
rect 114212 -480 114324 240
rect 115164 -480 115276 240
rect 116116 -480 116228 240
rect 117068 -480 117180 240
rect 118020 -480 118132 240
rect 118972 -480 119084 240
rect 119924 -480 120036 240
rect 120876 -480 120988 240
rect 121828 -480 121940 240
rect 122780 -480 122892 240
rect 123732 -480 123844 240
rect 124684 -480 124796 240
rect 125636 -480 125748 240
rect 126588 -480 126700 240
rect 127540 -480 127652 240
rect 128492 -480 128604 240
rect 129444 -480 129556 240
rect 130396 -480 130508 240
rect 131348 -480 131460 240
rect 132300 -480 132412 240
rect 133252 -480 133364 240
rect 134204 -480 134316 240
rect 135156 -480 135268 240
rect 136108 -480 136220 240
rect 137060 -480 137172 240
rect 138012 -480 138124 240
rect 138964 -480 139076 240
rect 139916 -480 140028 240
rect 140868 -480 140980 240
rect 141820 -480 141932 240
rect 142772 -480 142884 240
rect 143724 -480 143836 240
rect 144676 -480 144788 240
rect 145628 -480 145740 240
rect 146580 -480 146692 240
rect 147532 -480 147644 240
rect 148484 -480 148596 240
rect 149436 -480 149548 240
rect 150388 -480 150500 240
rect 151340 -480 151452 240
rect 152292 -480 152404 240
rect 153244 -480 153356 240
rect 154196 -480 154308 240
rect 155148 -480 155260 240
rect 156100 -480 156212 240
rect 157052 -480 157164 240
rect 158004 -480 158116 240
rect 158956 -480 159068 240
rect 159908 -480 160020 240
rect 160860 -480 160972 240
rect 161812 -480 161924 240
rect 162764 -480 162876 240
rect 163716 -480 163828 240
rect 164668 -480 164780 240
rect 165620 -480 165732 240
rect 166572 -480 166684 240
rect 167524 -480 167636 240
rect 168476 -480 168588 240
rect 169428 -480 169540 240
rect 170380 -480 170492 240
rect 171332 -480 171444 240
rect 172284 -480 172396 240
rect 173236 -480 173348 240
rect 174188 -480 174300 240
rect 175140 -480 175252 240
rect 176092 -480 176204 240
rect 177044 -480 177156 240
rect 177996 -480 178108 240
rect 178948 -480 179060 240
rect 179900 -480 180012 240
rect 180852 -480 180964 240
rect 181804 -480 181916 240
rect 182756 -480 182868 240
rect 183708 -480 183820 240
rect 184660 -480 184772 240
rect 185612 -480 185724 240
rect 186564 -480 186676 240
rect 187516 -480 187628 240
rect 188468 -480 188580 240
rect 189420 -480 189532 240
rect 190372 -480 190484 240
rect 191324 -480 191436 240
rect 192276 -480 192388 240
rect 193228 -480 193340 240
rect 194180 -480 194292 240
rect 195132 -480 195244 240
rect 196084 -480 196196 240
rect 197036 -480 197148 240
rect 197988 -480 198100 240
rect 198940 -480 199052 240
rect 199892 -480 200004 240
rect 200844 -480 200956 240
rect 201796 -480 201908 240
rect 202748 -480 202860 240
rect 203700 -480 203812 240
rect 204652 -480 204764 240
rect 205604 -480 205716 240
rect 206556 -480 206668 240
rect 207508 -480 207620 240
rect 208460 -480 208572 240
rect 209412 -480 209524 240
rect 210364 -480 210476 240
rect 211316 -480 211428 240
rect 212268 -480 212380 240
rect 213220 -480 213332 240
rect 214172 -480 214284 240
rect 215124 -480 215236 240
rect 216076 -480 216188 240
rect 217028 -480 217140 240
rect 217980 -480 218092 240
rect 218932 -480 219044 240
rect 219884 -480 219996 240
rect 220836 -480 220948 240
rect 221788 -480 221900 240
rect 222740 -480 222852 240
rect 223692 -480 223804 240
rect 224644 -480 224756 240
rect 225596 -480 225708 240
rect 226548 -480 226660 240
rect 227500 -480 227612 240
rect 228452 -480 228564 240
rect 229404 -480 229516 240
rect 230356 -480 230468 240
rect 231308 -480 231420 240
rect 232260 -480 232372 240
rect 233212 -480 233324 240
rect 234164 -480 234276 240
rect 235116 -480 235228 240
rect 236068 -480 236180 240
rect 237020 -480 237132 240
rect 237972 -480 238084 240
rect 238924 -480 239036 240
rect 239876 -480 239988 240
rect 240828 -480 240940 240
rect 241780 -480 241892 240
rect 242732 -480 242844 240
rect 243684 -480 243796 240
rect 244636 -480 244748 240
rect 245588 -480 245700 240
rect 246540 -480 246652 240
rect 247492 -480 247604 240
rect 248444 -480 248556 240
rect 249396 -480 249508 240
rect 250348 -480 250460 240
rect 251300 -480 251412 240
rect 252252 -480 252364 240
rect 253204 -480 253316 240
rect 254156 -480 254268 240
rect 255108 -480 255220 240
rect 256060 -480 256172 240
rect 257012 -480 257124 240
rect 257964 -480 258076 240
rect 258916 -480 259028 240
rect 259868 -480 259980 240
rect 260820 -480 260932 240
rect 261772 -480 261884 240
rect 262724 -480 262836 240
rect 263676 -480 263788 240
rect 264628 -480 264740 240
rect 265580 -480 265692 240
rect 266532 -480 266644 240
rect 267484 -480 267596 240
rect 268436 -480 268548 240
rect 269388 -480 269500 240
rect 270340 -480 270452 240
rect 271292 -480 271404 240
rect 272244 -480 272356 240
rect 273196 -480 273308 240
rect 274148 -480 274260 240
rect 275100 -480 275212 240
rect 276052 -480 276164 240
rect 277004 -480 277116 240
rect 277956 -480 278068 240
rect 278908 -480 279020 240
rect 279860 -480 279972 240
rect 280812 -480 280924 240
rect 281764 -480 281876 240
rect 282716 -480 282828 240
rect 283668 -480 283780 240
rect 284620 -480 284732 240
rect 285572 -480 285684 240
rect 286524 -480 286636 240
rect 287476 -480 287588 240
rect 288428 -480 288540 240
rect 289380 -480 289492 240
rect 290332 -480 290444 240
rect 291284 -480 291396 240
rect 292236 -480 292348 240
<< obsm2 >>
rect 2086 297750 5486 297850
rect 5658 297750 16518 297850
rect 16690 297750 27550 297850
rect 27722 297750 38582 297850
rect 38754 297750 49614 297850
rect 49786 297750 60646 297850
rect 60818 297750 71678 297850
rect 71850 297750 82710 297850
rect 82882 297750 93742 297850
rect 93914 297750 104774 297850
rect 104946 297750 115806 297850
rect 115978 297750 126838 297850
rect 127010 297750 137870 297850
rect 138042 297750 148902 297850
rect 149074 297750 159934 297850
rect 160106 297750 170966 297850
rect 171138 297750 181998 297850
rect 182170 297750 193030 297850
rect 193202 297750 204062 297850
rect 204234 297750 215094 297850
rect 215266 297750 226126 297850
rect 226298 297750 237158 297850
rect 237330 297750 248190 297850
rect 248362 297750 259222 297850
rect 259394 297750 270254 297850
rect 270426 297750 281286 297850
rect 281458 297750 292318 297850
rect 292490 297750 297178 297850
rect 2086 270 297178 297750
rect 2086 196 5654 270
rect 5826 196 6606 270
rect 6778 196 7558 270
rect 7730 196 8510 270
rect 8682 196 9462 270
rect 9634 196 10414 270
rect 10586 196 11366 270
rect 11538 196 12318 270
rect 12490 196 13270 270
rect 13442 196 14222 270
rect 14394 196 15174 270
rect 15346 196 16126 270
rect 16298 196 17078 270
rect 17250 196 18030 270
rect 18202 196 18982 270
rect 19154 196 19934 270
rect 20106 196 20886 270
rect 21058 196 21838 270
rect 22010 196 22790 270
rect 22962 196 23742 270
rect 23914 196 24694 270
rect 24866 196 25646 270
rect 25818 196 26598 270
rect 26770 196 27550 270
rect 27722 196 28502 270
rect 28674 196 29454 270
rect 29626 196 30406 270
rect 30578 196 31358 270
rect 31530 196 32310 270
rect 32482 196 33262 270
rect 33434 196 34214 270
rect 34386 196 35166 270
rect 35338 196 36118 270
rect 36290 196 37070 270
rect 37242 196 38022 270
rect 38194 196 38974 270
rect 39146 196 39926 270
rect 40098 196 40878 270
rect 41050 196 41830 270
rect 42002 196 42782 270
rect 42954 196 43734 270
rect 43906 196 44686 270
rect 44858 196 45638 270
rect 45810 196 46590 270
rect 46762 196 47542 270
rect 47714 196 48494 270
rect 48666 196 49446 270
rect 49618 196 50398 270
rect 50570 196 51350 270
rect 51522 196 52302 270
rect 52474 196 53254 270
rect 53426 196 54206 270
rect 54378 196 55158 270
rect 55330 196 56110 270
rect 56282 196 57062 270
rect 57234 196 58014 270
rect 58186 196 58966 270
rect 59138 196 59918 270
rect 60090 196 60870 270
rect 61042 196 61822 270
rect 61994 196 62774 270
rect 62946 196 63726 270
rect 63898 196 64678 270
rect 64850 196 65630 270
rect 65802 196 66582 270
rect 66754 196 67534 270
rect 67706 196 68486 270
rect 68658 196 69438 270
rect 69610 196 70390 270
rect 70562 196 71342 270
rect 71514 196 72294 270
rect 72466 196 73246 270
rect 73418 196 74198 270
rect 74370 196 75150 270
rect 75322 196 76102 270
rect 76274 196 77054 270
rect 77226 196 78006 270
rect 78178 196 78958 270
rect 79130 196 79910 270
rect 80082 196 80862 270
rect 81034 196 81814 270
rect 81986 196 82766 270
rect 82938 196 83718 270
rect 83890 196 84670 270
rect 84842 196 85622 270
rect 85794 196 86574 270
rect 86746 196 87526 270
rect 87698 196 88478 270
rect 88650 196 89430 270
rect 89602 196 90382 270
rect 90554 196 91334 270
rect 91506 196 92286 270
rect 92458 196 93238 270
rect 93410 196 94190 270
rect 94362 196 95142 270
rect 95314 196 96094 270
rect 96266 196 97046 270
rect 97218 196 97998 270
rect 98170 196 98950 270
rect 99122 196 99902 270
rect 100074 196 100854 270
rect 101026 196 101806 270
rect 101978 196 102758 270
rect 102930 196 103710 270
rect 103882 196 104662 270
rect 104834 196 105614 270
rect 105786 196 106566 270
rect 106738 196 107518 270
rect 107690 196 108470 270
rect 108642 196 109422 270
rect 109594 196 110374 270
rect 110546 196 111326 270
rect 111498 196 112278 270
rect 112450 196 113230 270
rect 113402 196 114182 270
rect 114354 196 115134 270
rect 115306 196 116086 270
rect 116258 196 117038 270
rect 117210 196 117990 270
rect 118162 196 118942 270
rect 119114 196 119894 270
rect 120066 196 120846 270
rect 121018 196 121798 270
rect 121970 196 122750 270
rect 122922 196 123702 270
rect 123874 196 124654 270
rect 124826 196 125606 270
rect 125778 196 126558 270
rect 126730 196 127510 270
rect 127682 196 128462 270
rect 128634 196 129414 270
rect 129586 196 130366 270
rect 130538 196 131318 270
rect 131490 196 132270 270
rect 132442 196 133222 270
rect 133394 196 134174 270
rect 134346 196 135126 270
rect 135298 196 136078 270
rect 136250 196 137030 270
rect 137202 196 137982 270
rect 138154 196 138934 270
rect 139106 196 139886 270
rect 140058 196 140838 270
rect 141010 196 141790 270
rect 141962 196 142742 270
rect 142914 196 143694 270
rect 143866 196 144646 270
rect 144818 196 145598 270
rect 145770 196 146550 270
rect 146722 196 147502 270
rect 147674 196 148454 270
rect 148626 196 149406 270
rect 149578 196 150358 270
rect 150530 196 151310 270
rect 151482 196 152262 270
rect 152434 196 153214 270
rect 153386 196 154166 270
rect 154338 196 155118 270
rect 155290 196 156070 270
rect 156242 196 157022 270
rect 157194 196 157974 270
rect 158146 196 158926 270
rect 159098 196 159878 270
rect 160050 196 160830 270
rect 161002 196 161782 270
rect 161954 196 162734 270
rect 162906 196 163686 270
rect 163858 196 164638 270
rect 164810 196 165590 270
rect 165762 196 166542 270
rect 166714 196 167494 270
rect 167666 196 168446 270
rect 168618 196 169398 270
rect 169570 196 170350 270
rect 170522 196 171302 270
rect 171474 196 172254 270
rect 172426 196 173206 270
rect 173378 196 174158 270
rect 174330 196 175110 270
rect 175282 196 176062 270
rect 176234 196 177014 270
rect 177186 196 177966 270
rect 178138 196 178918 270
rect 179090 196 179870 270
rect 180042 196 180822 270
rect 180994 196 181774 270
rect 181946 196 182726 270
rect 182898 196 183678 270
rect 183850 196 184630 270
rect 184802 196 185582 270
rect 185754 196 186534 270
rect 186706 196 187486 270
rect 187658 196 188438 270
rect 188610 196 189390 270
rect 189562 196 190342 270
rect 190514 196 191294 270
rect 191466 196 192246 270
rect 192418 196 193198 270
rect 193370 196 194150 270
rect 194322 196 195102 270
rect 195274 196 196054 270
rect 196226 196 197006 270
rect 197178 196 197958 270
rect 198130 196 198910 270
rect 199082 196 199862 270
rect 200034 196 200814 270
rect 200986 196 201766 270
rect 201938 196 202718 270
rect 202890 196 203670 270
rect 203842 196 204622 270
rect 204794 196 205574 270
rect 205746 196 206526 270
rect 206698 196 207478 270
rect 207650 196 208430 270
rect 208602 196 209382 270
rect 209554 196 210334 270
rect 210506 196 211286 270
rect 211458 196 212238 270
rect 212410 196 213190 270
rect 213362 196 214142 270
rect 214314 196 215094 270
rect 215266 196 216046 270
rect 216218 196 216998 270
rect 217170 196 217950 270
rect 218122 196 218902 270
rect 219074 196 219854 270
rect 220026 196 220806 270
rect 220978 196 221758 270
rect 221930 196 222710 270
rect 222882 196 223662 270
rect 223834 196 224614 270
rect 224786 196 225566 270
rect 225738 196 226518 270
rect 226690 196 227470 270
rect 227642 196 228422 270
rect 228594 196 229374 270
rect 229546 196 230326 270
rect 230498 196 231278 270
rect 231450 196 232230 270
rect 232402 196 233182 270
rect 233354 196 234134 270
rect 234306 196 235086 270
rect 235258 196 236038 270
rect 236210 196 236990 270
rect 237162 196 237942 270
rect 238114 196 238894 270
rect 239066 196 239846 270
rect 240018 196 240798 270
rect 240970 196 241750 270
rect 241922 196 242702 270
rect 242874 196 243654 270
rect 243826 196 244606 270
rect 244778 196 245558 270
rect 245730 196 246510 270
rect 246682 196 247462 270
rect 247634 196 248414 270
rect 248586 196 249366 270
rect 249538 196 250318 270
rect 250490 196 251270 270
rect 251442 196 252222 270
rect 252394 196 253174 270
rect 253346 196 254126 270
rect 254298 196 255078 270
rect 255250 196 256030 270
rect 256202 196 256982 270
rect 257154 196 257934 270
rect 258106 196 258886 270
rect 259058 196 259838 270
rect 260010 196 260790 270
rect 260962 196 261742 270
rect 261914 196 262694 270
rect 262866 196 263646 270
rect 263818 196 264598 270
rect 264770 196 265550 270
rect 265722 196 266502 270
rect 266674 196 267454 270
rect 267626 196 268406 270
rect 268578 196 269358 270
rect 269530 196 270310 270
rect 270482 196 271262 270
rect 271434 196 272214 270
rect 272386 196 273166 270
rect 273338 196 274118 270
rect 274290 196 275070 270
rect 275242 196 276022 270
rect 276194 196 276974 270
rect 277146 196 277926 270
rect 278098 196 278878 270
rect 279050 196 279830 270
rect 280002 196 280782 270
rect 280954 196 281734 270
rect 281906 196 282686 270
rect 282858 196 283638 270
rect 283810 196 284590 270
rect 284762 196 285542 270
rect 285714 196 286494 270
rect 286666 196 287446 270
rect 287618 196 288398 270
rect 288570 196 289350 270
rect 289522 196 290302 270
rect 290474 196 291254 270
rect 291426 196 292206 270
rect 292378 196 297178 270
<< metal3 >>
rect 297780 294308 298500 294420
rect -480 293580 240 293692
rect 297780 287700 298500 287812
rect -480 286524 240 286636
rect 297780 281092 298500 281204
rect -480 279468 240 279580
rect 297780 274484 298500 274596
rect -480 272412 240 272524
rect 297780 267876 298500 267988
rect -480 265356 240 265468
rect 297780 261268 298500 261380
rect -480 258300 240 258412
rect 297780 254660 298500 254772
rect -480 251244 240 251356
rect 297780 248052 298500 248164
rect -480 244188 240 244300
rect 297780 241444 298500 241556
rect -480 237132 240 237244
rect 297780 234836 298500 234948
rect -480 230076 240 230188
rect 297780 228228 298500 228340
rect -480 223020 240 223132
rect 297780 221620 298500 221732
rect -480 215964 240 216076
rect 297780 215012 298500 215124
rect -480 208908 240 209020
rect 297780 208404 298500 208516
rect -480 201852 240 201964
rect 297780 201796 298500 201908
rect 297780 195188 298500 195300
rect -480 194796 240 194908
rect 297780 188580 298500 188692
rect -480 187740 240 187852
rect 297780 181972 298500 182084
rect -480 180684 240 180796
rect 297780 175364 298500 175476
rect -480 173628 240 173740
rect 297780 168756 298500 168868
rect -480 166572 240 166684
rect 297780 162148 298500 162260
rect -480 159516 240 159628
rect 297780 155540 298500 155652
rect -480 152460 240 152572
rect 297780 148932 298500 149044
rect -480 145404 240 145516
rect 297780 142324 298500 142436
rect -480 138348 240 138460
rect 297780 135716 298500 135828
rect -480 131292 240 131404
rect 297780 129108 298500 129220
rect -480 124236 240 124348
rect 297780 122500 298500 122612
rect -480 117180 240 117292
rect 297780 115892 298500 116004
rect -480 110124 240 110236
rect 297780 109284 298500 109396
rect -480 103068 240 103180
rect 297780 102676 298500 102788
rect -480 96012 240 96124
rect 297780 96068 298500 96180
rect 297780 89460 298500 89572
rect -480 88956 240 89068
rect 297780 82852 298500 82964
rect -480 81900 240 82012
rect 297780 76244 298500 76356
rect -480 74844 240 74956
rect 297780 69636 298500 69748
rect -480 67788 240 67900
rect 297780 63028 298500 63140
rect -480 60732 240 60844
rect 297780 56420 298500 56532
rect -480 53676 240 53788
rect 297780 49812 298500 49924
rect -480 46620 240 46732
rect 297780 43204 298500 43316
rect -480 39564 240 39676
rect 297780 36596 298500 36708
rect -480 32508 240 32620
rect 297780 29988 298500 30100
rect -480 25452 240 25564
rect 297780 23380 298500 23492
rect -480 18396 240 18508
rect 297780 16772 298500 16884
rect -480 11340 240 11452
rect 297780 10164 298500 10276
rect -480 4284 240 4396
rect 297780 3556 298500 3668
<< obsm3 >>
rect 182 294450 297850 295666
rect 182 294278 297750 294450
rect 182 293722 297850 294278
rect 270 293550 297850 293722
rect 182 287842 297850 293550
rect 182 287670 297750 287842
rect 182 286666 297850 287670
rect 270 286494 297850 286666
rect 182 281234 297850 286494
rect 182 281062 297750 281234
rect 182 279610 297850 281062
rect 270 279438 297850 279610
rect 182 274626 297850 279438
rect 182 274454 297750 274626
rect 182 272554 297850 274454
rect 270 272382 297850 272554
rect 182 268018 297850 272382
rect 182 267846 297750 268018
rect 182 265498 297850 267846
rect 270 265326 297850 265498
rect 182 261410 297850 265326
rect 182 261238 297750 261410
rect 182 258442 297850 261238
rect 270 258270 297850 258442
rect 182 254802 297850 258270
rect 182 254630 297750 254802
rect 182 251386 297850 254630
rect 270 251214 297850 251386
rect 182 248194 297850 251214
rect 182 248022 297750 248194
rect 182 244330 297850 248022
rect 270 244158 297850 244330
rect 182 241586 297850 244158
rect 182 241414 297750 241586
rect 182 237274 297850 241414
rect 270 237102 297850 237274
rect 182 234978 297850 237102
rect 182 234806 297750 234978
rect 182 230218 297850 234806
rect 270 230046 297850 230218
rect 182 228370 297850 230046
rect 182 228198 297750 228370
rect 182 223162 297850 228198
rect 270 222990 297850 223162
rect 182 221762 297850 222990
rect 182 221590 297750 221762
rect 182 216106 297850 221590
rect 270 215934 297850 216106
rect 182 215154 297850 215934
rect 182 214982 297750 215154
rect 182 209050 297850 214982
rect 270 208878 297850 209050
rect 182 208546 297850 208878
rect 182 208374 297750 208546
rect 182 201994 297850 208374
rect 270 201938 297850 201994
rect 270 201822 297750 201938
rect 182 201766 297750 201822
rect 182 195330 297850 201766
rect 182 195158 297750 195330
rect 182 194938 297850 195158
rect 270 194766 297850 194938
rect 182 188722 297850 194766
rect 182 188550 297750 188722
rect 182 187882 297850 188550
rect 270 187710 297850 187882
rect 182 182114 297850 187710
rect 182 181942 297750 182114
rect 182 180826 297850 181942
rect 270 180654 297850 180826
rect 182 175506 297850 180654
rect 182 175334 297750 175506
rect 182 173770 297850 175334
rect 270 173598 297850 173770
rect 182 168898 297850 173598
rect 182 168726 297750 168898
rect 182 166714 297850 168726
rect 270 166542 297850 166714
rect 182 162290 297850 166542
rect 182 162118 297750 162290
rect 182 159658 297850 162118
rect 270 159486 297850 159658
rect 182 155682 297850 159486
rect 182 155510 297750 155682
rect 182 152602 297850 155510
rect 270 152430 297850 152602
rect 182 149074 297850 152430
rect 182 148902 297750 149074
rect 182 145546 297850 148902
rect 270 145374 297850 145546
rect 182 142466 297850 145374
rect 182 142294 297750 142466
rect 182 138490 297850 142294
rect 270 138318 297850 138490
rect 182 135858 297850 138318
rect 182 135686 297750 135858
rect 182 131434 297850 135686
rect 270 131262 297850 131434
rect 182 129250 297850 131262
rect 182 129078 297750 129250
rect 182 124378 297850 129078
rect 270 124206 297850 124378
rect 182 122642 297850 124206
rect 182 122470 297750 122642
rect 182 117322 297850 122470
rect 270 117150 297850 117322
rect 182 116034 297850 117150
rect 182 115862 297750 116034
rect 182 110266 297850 115862
rect 270 110094 297850 110266
rect 182 109426 297850 110094
rect 182 109254 297750 109426
rect 182 103210 297850 109254
rect 270 103038 297850 103210
rect 182 102818 297850 103038
rect 182 102646 297750 102818
rect 182 96210 297850 102646
rect 182 96154 297750 96210
rect 270 96038 297750 96154
rect 270 95982 297850 96038
rect 182 89602 297850 95982
rect 182 89430 297750 89602
rect 182 89098 297850 89430
rect 270 88926 297850 89098
rect 182 82994 297850 88926
rect 182 82822 297750 82994
rect 182 82042 297850 82822
rect 270 81870 297850 82042
rect 182 76386 297850 81870
rect 182 76214 297750 76386
rect 182 74986 297850 76214
rect 270 74814 297850 74986
rect 182 69778 297850 74814
rect 182 69606 297750 69778
rect 182 67930 297850 69606
rect 270 67758 297850 67930
rect 182 63170 297850 67758
rect 182 62998 297750 63170
rect 182 60874 297850 62998
rect 270 60702 297850 60874
rect 182 56562 297850 60702
rect 182 56390 297750 56562
rect 182 53818 297850 56390
rect 270 53646 297850 53818
rect 182 49954 297850 53646
rect 182 49782 297750 49954
rect 182 46762 297850 49782
rect 270 46590 297850 46762
rect 182 43346 297850 46590
rect 182 43174 297750 43346
rect 182 39706 297850 43174
rect 270 39534 297850 39706
rect 182 36738 297850 39534
rect 182 36566 297750 36738
rect 182 32650 297850 36566
rect 270 32478 297850 32650
rect 182 30130 297850 32478
rect 182 29958 297750 30130
rect 182 25594 297850 29958
rect 270 25422 297850 25594
rect 182 23522 297850 25422
rect 182 23350 297750 23522
rect 182 18538 297850 23350
rect 270 18366 297850 18538
rect 182 16914 297850 18366
rect 182 16742 297750 16914
rect 182 11482 297850 16742
rect 270 11310 297850 11482
rect 182 10306 297850 11310
rect 182 10134 297750 10306
rect 182 4426 297850 10134
rect 270 4254 297850 4426
rect 182 3698 297850 4254
rect 182 3526 297750 3698
rect 182 2086 297850 3526
<< metal4 >>
rect -958 -822 -648 299134
rect -478 -342 -168 298654
rect 1577 -822 1887 299134
rect 3437 -822 3747 299134
rect 10577 -822 10887 299134
rect 12437 -822 12747 299134
rect 19577 -822 19887 299134
rect 21437 -822 21747 299134
rect 28577 -822 28887 299134
rect 30437 -822 30747 299134
rect 37577 -822 37887 299134
rect 39437 -822 39747 299134
rect 46577 -822 46887 299134
rect 48437 -822 48747 299134
rect 55577 -822 55887 299134
rect 57437 -822 57747 299134
rect 64577 -822 64887 299134
rect 66437 -822 66747 299134
rect 73577 -822 73887 299134
rect 75437 -822 75747 299134
rect 82577 -822 82887 299134
rect 84437 -822 84747 299134
rect 91577 -822 91887 299134
rect 93437 -822 93747 299134
rect 100577 -822 100887 299134
rect 102437 -822 102747 299134
rect 109577 -822 109887 299134
rect 111437 -822 111747 299134
rect 118577 229771 118887 299134
rect 120437 229771 120747 299134
rect 127577 229771 127887 299134
rect 129437 229771 129747 299134
rect 136577 229771 136887 299134
rect 138437 229771 138747 299134
rect 145577 229771 145887 299134
rect 147437 229771 147747 299134
rect 154577 229771 154887 299134
rect 156437 229771 156747 299134
rect 163577 229771 163887 299134
rect 165437 229771 165747 299134
rect 172577 229771 172887 299134
rect 174437 229771 174747 299134
rect 181577 229771 181887 299134
rect 183437 229771 183747 299134
rect 190577 229771 190887 299134
rect 192437 229771 192747 299134
rect 199577 229771 199887 299134
rect 201437 229771 201747 299134
rect 118577 -822 118887 168709
rect 120437 -822 120747 168709
rect 127577 -822 127887 168709
rect 129437 -822 129747 168709
rect 136577 -822 136887 168709
rect 138437 -822 138747 168709
rect 145577 -822 145887 168709
rect 147437 -822 147747 168709
rect 154577 -822 154887 168709
rect 156437 -822 156747 168709
rect 163577 -822 163887 168709
rect 165437 -822 165747 168709
rect 172577 -822 172887 168709
rect 174437 -822 174747 168709
rect 181577 -822 181887 168709
rect 183437 -822 183747 168709
rect 190577 -822 190887 168709
rect 192437 -822 192747 168709
rect 199577 -822 199887 168709
rect 201437 -822 201747 168709
rect 208577 -822 208887 299134
rect 210437 -822 210747 299134
rect 217577 -822 217887 299134
rect 219437 -822 219747 299134
rect 226577 -822 226887 299134
rect 228437 -822 228747 299134
rect 235577 -822 235887 299134
rect 237437 -822 237747 299134
rect 244577 -822 244887 299134
rect 246437 -822 246747 299134
rect 253577 -822 253887 299134
rect 255437 -822 255747 299134
rect 262577 -822 262887 299134
rect 264437 -822 264747 299134
rect 271577 -822 271887 299134
rect 273437 -822 273747 299134
rect 280577 -822 280887 299134
rect 282437 -822 282747 299134
rect 289577 -822 289887 299134
rect 291437 -822 291747 299134
rect 298200 -342 298510 298654
rect 298680 -822 298990 299134
<< obsm4 >>
rect 119250 169737 205126 228743
<< metal5 >>
rect -958 298824 298990 299134
rect -478 298344 298510 298654
rect -958 292913 298990 293223
rect -958 289913 298990 290223
rect -958 283913 298990 284223
rect -958 280913 298990 281223
rect -958 274913 298990 275223
rect -958 271913 298990 272223
rect -958 265913 298990 266223
rect -958 262913 298990 263223
rect -958 256913 298990 257223
rect -958 253913 298990 254223
rect -958 247913 298990 248223
rect -958 244913 298990 245223
rect -958 238913 298990 239223
rect -958 235913 298990 236223
rect -958 229913 298990 230223
rect -958 226913 298990 227223
rect -958 220913 298990 221223
rect -958 217913 298990 218223
rect -958 211913 298990 212223
rect -958 208913 298990 209223
rect -958 202913 298990 203223
rect -958 199913 298990 200223
rect -958 193913 298990 194223
rect -958 190913 298990 191223
rect -958 184913 298990 185223
rect -958 181913 298990 182223
rect -958 175913 298990 176223
rect -958 172913 298990 173223
rect -958 166913 298990 167223
rect -958 163913 298990 164223
rect -958 157913 298990 158223
rect -958 154913 298990 155223
rect -958 148913 298990 149223
rect -958 145913 298990 146223
rect -958 139913 298990 140223
rect -958 136913 298990 137223
rect -958 130913 298990 131223
rect -958 127913 298990 128223
rect -958 121913 298990 122223
rect -958 118913 298990 119223
rect -958 112913 298990 113223
rect -958 109913 298990 110223
rect -958 103913 298990 104223
rect -958 100913 298990 101223
rect -958 94913 298990 95223
rect -958 91913 298990 92223
rect -958 85913 298990 86223
rect -958 82913 298990 83223
rect -958 76913 298990 77223
rect -958 73913 298990 74223
rect -958 67913 298990 68223
rect -958 64913 298990 65223
rect -958 58913 298990 59223
rect -958 55913 298990 56223
rect -958 49913 298990 50223
rect -958 46913 298990 47223
rect -958 40913 298990 41223
rect -958 37913 298990 38223
rect -958 31913 298990 32223
rect -958 28913 298990 29223
rect -958 22913 298990 23223
rect -958 19913 298990 20223
rect -958 13913 298990 14223
rect -958 10913 298990 11223
rect -958 4913 298990 5223
rect -958 1913 298990 2223
rect -478 -342 298510 -32
rect -958 -822 298990 -512
<< labels >>
rlabel metal3 s 297780 3556 298500 3668 6 io_in[0]
port 1 nsew signal input
rlabel metal3 s 297780 201796 298500 201908 6 io_in[10]
port 2 nsew signal input
rlabel metal3 s 297780 221620 298500 221732 6 io_in[11]
port 3 nsew signal input
rlabel metal3 s 297780 241444 298500 241556 6 io_in[12]
port 4 nsew signal input
rlabel metal3 s 297780 261268 298500 261380 6 io_in[13]
port 5 nsew signal input
rlabel metal3 s 297780 281092 298500 281204 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 292348 297780 292460 298500 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 259252 297780 259364 298500 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 226156 297780 226268 298500 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 193060 297780 193172 298500 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 159964 297780 160076 298500 6 io_in[19]
port 11 nsew signal input
rlabel metal3 s 297780 23380 298500 23492 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 126868 297780 126980 298500 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 93772 297780 93884 298500 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 60676 297780 60788 298500 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 27580 297780 27692 298500 6 io_in[23]
port 16 nsew signal input
rlabel metal3 s -480 293580 240 293692 4 io_in[24]
port 17 nsew signal input
rlabel metal3 s -480 272412 240 272524 4 io_in[25]
port 18 nsew signal input
rlabel metal3 s -480 251244 240 251356 4 io_in[26]
port 19 nsew signal input
rlabel metal3 s -480 230076 240 230188 4 io_in[27]
port 20 nsew signal input
rlabel metal3 s -480 208908 240 209020 4 io_in[28]
port 21 nsew signal input
rlabel metal3 s -480 187740 240 187852 4 io_in[29]
port 22 nsew signal input
rlabel metal3 s 297780 43204 298500 43316 6 io_in[2]
port 23 nsew signal input
rlabel metal3 s -480 166572 240 166684 4 io_in[30]
port 24 nsew signal input
rlabel metal3 s -480 145404 240 145516 4 io_in[31]
port 25 nsew signal input
rlabel metal3 s -480 124236 240 124348 4 io_in[32]
port 26 nsew signal input
rlabel metal3 s -480 103068 240 103180 4 io_in[33]
port 27 nsew signal input
rlabel metal3 s -480 81900 240 82012 4 io_in[34]
port 28 nsew signal input
rlabel metal3 s -480 60732 240 60844 4 io_in[35]
port 29 nsew signal input
rlabel metal3 s -480 39564 240 39676 4 io_in[36]
port 30 nsew signal input
rlabel metal3 s -480 18396 240 18508 4 io_in[37]
port 31 nsew signal input
rlabel metal3 s 297780 63028 298500 63140 6 io_in[3]
port 32 nsew signal input
rlabel metal3 s 297780 82852 298500 82964 6 io_in[4]
port 33 nsew signal input
rlabel metal3 s 297780 102676 298500 102788 6 io_in[5]
port 34 nsew signal input
rlabel metal3 s 297780 122500 298500 122612 6 io_in[6]
port 35 nsew signal input
rlabel metal3 s 297780 142324 298500 142436 6 io_in[7]
port 36 nsew signal input
rlabel metal3 s 297780 162148 298500 162260 6 io_in[8]
port 37 nsew signal input
rlabel metal3 s 297780 181972 298500 182084 6 io_in[9]
port 38 nsew signal input
rlabel metal3 s 297780 16772 298500 16884 6 io_oeb[0]
port 39 nsew signal output
rlabel metal3 s 297780 215012 298500 215124 6 io_oeb[10]
port 40 nsew signal output
rlabel metal3 s 297780 234836 298500 234948 6 io_oeb[11]
port 41 nsew signal output
rlabel metal3 s 297780 254660 298500 254772 6 io_oeb[12]
port 42 nsew signal output
rlabel metal3 s 297780 274484 298500 274596 6 io_oeb[13]
port 43 nsew signal output
rlabel metal3 s 297780 294308 298500 294420 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 270284 297780 270396 298500 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 237188 297780 237300 298500 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 204092 297780 204204 298500 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 170996 297780 171108 298500 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 137900 297780 138012 298500 6 io_oeb[19]
port 49 nsew signal output
rlabel metal3 s 297780 36596 298500 36708 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 104804 297780 104916 298500 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 71708 297780 71820 298500 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 38612 297780 38724 298500 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 5516 297780 5628 298500 6 io_oeb[23]
port 54 nsew signal output
rlabel metal3 s -480 279468 240 279580 4 io_oeb[24]
port 55 nsew signal output
rlabel metal3 s -480 258300 240 258412 4 io_oeb[25]
port 56 nsew signal output
rlabel metal3 s -480 237132 240 237244 4 io_oeb[26]
port 57 nsew signal output
rlabel metal3 s -480 215964 240 216076 4 io_oeb[27]
port 58 nsew signal output
rlabel metal3 s -480 194796 240 194908 4 io_oeb[28]
port 59 nsew signal output
rlabel metal3 s -480 173628 240 173740 4 io_oeb[29]
port 60 nsew signal output
rlabel metal3 s 297780 56420 298500 56532 6 io_oeb[2]
port 61 nsew signal output
rlabel metal3 s -480 152460 240 152572 4 io_oeb[30]
port 62 nsew signal output
rlabel metal3 s -480 131292 240 131404 4 io_oeb[31]
port 63 nsew signal output
rlabel metal3 s -480 110124 240 110236 4 io_oeb[32]
port 64 nsew signal output
rlabel metal3 s -480 88956 240 89068 4 io_oeb[33]
port 65 nsew signal output
rlabel metal3 s -480 67788 240 67900 4 io_oeb[34]
port 66 nsew signal output
rlabel metal3 s -480 46620 240 46732 4 io_oeb[35]
port 67 nsew signal output
rlabel metal3 s -480 25452 240 25564 4 io_oeb[36]
port 68 nsew signal output
rlabel metal3 s -480 4284 240 4396 4 io_oeb[37]
port 69 nsew signal output
rlabel metal3 s 297780 76244 298500 76356 6 io_oeb[3]
port 70 nsew signal output
rlabel metal3 s 297780 96068 298500 96180 6 io_oeb[4]
port 71 nsew signal output
rlabel metal3 s 297780 115892 298500 116004 6 io_oeb[5]
port 72 nsew signal output
rlabel metal3 s 297780 135716 298500 135828 6 io_oeb[6]
port 73 nsew signal output
rlabel metal3 s 297780 155540 298500 155652 6 io_oeb[7]
port 74 nsew signal output
rlabel metal3 s 297780 175364 298500 175476 6 io_oeb[8]
port 75 nsew signal output
rlabel metal3 s 297780 195188 298500 195300 6 io_oeb[9]
port 76 nsew signal output
rlabel metal3 s 297780 10164 298500 10276 6 io_out[0]
port 77 nsew signal output
rlabel metal3 s 297780 208404 298500 208516 6 io_out[10]
port 78 nsew signal output
rlabel metal3 s 297780 228228 298500 228340 6 io_out[11]
port 79 nsew signal output
rlabel metal3 s 297780 248052 298500 248164 6 io_out[12]
port 80 nsew signal output
rlabel metal3 s 297780 267876 298500 267988 6 io_out[13]
port 81 nsew signal output
rlabel metal3 s 297780 287700 298500 287812 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 281316 297780 281428 298500 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 248220 297780 248332 298500 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 215124 297780 215236 298500 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 182028 297780 182140 298500 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 148932 297780 149044 298500 6 io_out[19]
port 87 nsew signal output
rlabel metal3 s 297780 29988 298500 30100 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 115836 297780 115948 298500 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 82740 297780 82852 298500 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 49644 297780 49756 298500 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 16548 297780 16660 298500 6 io_out[23]
port 92 nsew signal output
rlabel metal3 s -480 286524 240 286636 4 io_out[24]
port 93 nsew signal output
rlabel metal3 s -480 265356 240 265468 4 io_out[25]
port 94 nsew signal output
rlabel metal3 s -480 244188 240 244300 4 io_out[26]
port 95 nsew signal output
rlabel metal3 s -480 223020 240 223132 4 io_out[27]
port 96 nsew signal output
rlabel metal3 s -480 201852 240 201964 4 io_out[28]
port 97 nsew signal output
rlabel metal3 s -480 180684 240 180796 4 io_out[29]
port 98 nsew signal output
rlabel metal3 s 297780 49812 298500 49924 6 io_out[2]
port 99 nsew signal output
rlabel metal3 s -480 159516 240 159628 4 io_out[30]
port 100 nsew signal output
rlabel metal3 s -480 138348 240 138460 4 io_out[31]
port 101 nsew signal output
rlabel metal3 s -480 117180 240 117292 4 io_out[32]
port 102 nsew signal output
rlabel metal3 s -480 96012 240 96124 4 io_out[33]
port 103 nsew signal output
rlabel metal3 s -480 74844 240 74956 4 io_out[34]
port 104 nsew signal output
rlabel metal3 s -480 53676 240 53788 4 io_out[35]
port 105 nsew signal output
rlabel metal3 s -480 32508 240 32620 4 io_out[36]
port 106 nsew signal output
rlabel metal3 s -480 11340 240 11452 4 io_out[37]
port 107 nsew signal output
rlabel metal3 s 297780 69636 298500 69748 6 io_out[3]
port 108 nsew signal output
rlabel metal3 s 297780 89460 298500 89572 6 io_out[4]
port 109 nsew signal output
rlabel metal3 s 297780 109284 298500 109396 6 io_out[5]
port 110 nsew signal output
rlabel metal3 s 297780 129108 298500 129220 6 io_out[6]
port 111 nsew signal output
rlabel metal3 s 297780 148932 298500 149044 6 io_out[7]
port 112 nsew signal output
rlabel metal3 s 297780 168756 298500 168868 6 io_out[8]
port 113 nsew signal output
rlabel metal3 s 297780 188580 298500 188692 6 io_out[9]
port 114 nsew signal output
rlabel metal2 s 106596 -480 106708 240 8 la_data_in[0]
port 115 nsew signal input
rlabel metal2 s 135156 -480 135268 240 8 la_data_in[10]
port 116 nsew signal input
rlabel metal2 s 138012 -480 138124 240 8 la_data_in[11]
port 117 nsew signal input
rlabel metal2 s 140868 -480 140980 240 8 la_data_in[12]
port 118 nsew signal input
rlabel metal2 s 143724 -480 143836 240 8 la_data_in[13]
port 119 nsew signal input
rlabel metal2 s 146580 -480 146692 240 8 la_data_in[14]
port 120 nsew signal input
rlabel metal2 s 149436 -480 149548 240 8 la_data_in[15]
port 121 nsew signal input
rlabel metal2 s 152292 -480 152404 240 8 la_data_in[16]
port 122 nsew signal input
rlabel metal2 s 155148 -480 155260 240 8 la_data_in[17]
port 123 nsew signal input
rlabel metal2 s 158004 -480 158116 240 8 la_data_in[18]
port 124 nsew signal input
rlabel metal2 s 160860 -480 160972 240 8 la_data_in[19]
port 125 nsew signal input
rlabel metal2 s 109452 -480 109564 240 8 la_data_in[1]
port 126 nsew signal input
rlabel metal2 s 163716 -480 163828 240 8 la_data_in[20]
port 127 nsew signal input
rlabel metal2 s 166572 -480 166684 240 8 la_data_in[21]
port 128 nsew signal input
rlabel metal2 s 169428 -480 169540 240 8 la_data_in[22]
port 129 nsew signal input
rlabel metal2 s 172284 -480 172396 240 8 la_data_in[23]
port 130 nsew signal input
rlabel metal2 s 175140 -480 175252 240 8 la_data_in[24]
port 131 nsew signal input
rlabel metal2 s 177996 -480 178108 240 8 la_data_in[25]
port 132 nsew signal input
rlabel metal2 s 180852 -480 180964 240 8 la_data_in[26]
port 133 nsew signal input
rlabel metal2 s 183708 -480 183820 240 8 la_data_in[27]
port 134 nsew signal input
rlabel metal2 s 186564 -480 186676 240 8 la_data_in[28]
port 135 nsew signal input
rlabel metal2 s 189420 -480 189532 240 8 la_data_in[29]
port 136 nsew signal input
rlabel metal2 s 112308 -480 112420 240 8 la_data_in[2]
port 137 nsew signal input
rlabel metal2 s 192276 -480 192388 240 8 la_data_in[30]
port 138 nsew signal input
rlabel metal2 s 195132 -480 195244 240 8 la_data_in[31]
port 139 nsew signal input
rlabel metal2 s 197988 -480 198100 240 8 la_data_in[32]
port 140 nsew signal input
rlabel metal2 s 200844 -480 200956 240 8 la_data_in[33]
port 141 nsew signal input
rlabel metal2 s 203700 -480 203812 240 8 la_data_in[34]
port 142 nsew signal input
rlabel metal2 s 206556 -480 206668 240 8 la_data_in[35]
port 143 nsew signal input
rlabel metal2 s 209412 -480 209524 240 8 la_data_in[36]
port 144 nsew signal input
rlabel metal2 s 212268 -480 212380 240 8 la_data_in[37]
port 145 nsew signal input
rlabel metal2 s 215124 -480 215236 240 8 la_data_in[38]
port 146 nsew signal input
rlabel metal2 s 217980 -480 218092 240 8 la_data_in[39]
port 147 nsew signal input
rlabel metal2 s 115164 -480 115276 240 8 la_data_in[3]
port 148 nsew signal input
rlabel metal2 s 220836 -480 220948 240 8 la_data_in[40]
port 149 nsew signal input
rlabel metal2 s 223692 -480 223804 240 8 la_data_in[41]
port 150 nsew signal input
rlabel metal2 s 226548 -480 226660 240 8 la_data_in[42]
port 151 nsew signal input
rlabel metal2 s 229404 -480 229516 240 8 la_data_in[43]
port 152 nsew signal input
rlabel metal2 s 232260 -480 232372 240 8 la_data_in[44]
port 153 nsew signal input
rlabel metal2 s 235116 -480 235228 240 8 la_data_in[45]
port 154 nsew signal input
rlabel metal2 s 237972 -480 238084 240 8 la_data_in[46]
port 155 nsew signal input
rlabel metal2 s 240828 -480 240940 240 8 la_data_in[47]
port 156 nsew signal input
rlabel metal2 s 243684 -480 243796 240 8 la_data_in[48]
port 157 nsew signal input
rlabel metal2 s 246540 -480 246652 240 8 la_data_in[49]
port 158 nsew signal input
rlabel metal2 s 118020 -480 118132 240 8 la_data_in[4]
port 159 nsew signal input
rlabel metal2 s 249396 -480 249508 240 8 la_data_in[50]
port 160 nsew signal input
rlabel metal2 s 252252 -480 252364 240 8 la_data_in[51]
port 161 nsew signal input
rlabel metal2 s 255108 -480 255220 240 8 la_data_in[52]
port 162 nsew signal input
rlabel metal2 s 257964 -480 258076 240 8 la_data_in[53]
port 163 nsew signal input
rlabel metal2 s 260820 -480 260932 240 8 la_data_in[54]
port 164 nsew signal input
rlabel metal2 s 263676 -480 263788 240 8 la_data_in[55]
port 165 nsew signal input
rlabel metal2 s 266532 -480 266644 240 8 la_data_in[56]
port 166 nsew signal input
rlabel metal2 s 269388 -480 269500 240 8 la_data_in[57]
port 167 nsew signal input
rlabel metal2 s 272244 -480 272356 240 8 la_data_in[58]
port 168 nsew signal input
rlabel metal2 s 275100 -480 275212 240 8 la_data_in[59]
port 169 nsew signal input
rlabel metal2 s 120876 -480 120988 240 8 la_data_in[5]
port 170 nsew signal input
rlabel metal2 s 277956 -480 278068 240 8 la_data_in[60]
port 171 nsew signal input
rlabel metal2 s 280812 -480 280924 240 8 la_data_in[61]
port 172 nsew signal input
rlabel metal2 s 283668 -480 283780 240 8 la_data_in[62]
port 173 nsew signal input
rlabel metal2 s 286524 -480 286636 240 8 la_data_in[63]
port 174 nsew signal input
rlabel metal2 s 123732 -480 123844 240 8 la_data_in[6]
port 175 nsew signal input
rlabel metal2 s 126588 -480 126700 240 8 la_data_in[7]
port 176 nsew signal input
rlabel metal2 s 129444 -480 129556 240 8 la_data_in[8]
port 177 nsew signal input
rlabel metal2 s 132300 -480 132412 240 8 la_data_in[9]
port 178 nsew signal input
rlabel metal2 s 107548 -480 107660 240 8 la_data_out[0]
port 179 nsew signal output
rlabel metal2 s 136108 -480 136220 240 8 la_data_out[10]
port 180 nsew signal output
rlabel metal2 s 138964 -480 139076 240 8 la_data_out[11]
port 181 nsew signal output
rlabel metal2 s 141820 -480 141932 240 8 la_data_out[12]
port 182 nsew signal output
rlabel metal2 s 144676 -480 144788 240 8 la_data_out[13]
port 183 nsew signal output
rlabel metal2 s 147532 -480 147644 240 8 la_data_out[14]
port 184 nsew signal output
rlabel metal2 s 150388 -480 150500 240 8 la_data_out[15]
port 185 nsew signal output
rlabel metal2 s 153244 -480 153356 240 8 la_data_out[16]
port 186 nsew signal output
rlabel metal2 s 156100 -480 156212 240 8 la_data_out[17]
port 187 nsew signal output
rlabel metal2 s 158956 -480 159068 240 8 la_data_out[18]
port 188 nsew signal output
rlabel metal2 s 161812 -480 161924 240 8 la_data_out[19]
port 189 nsew signal output
rlabel metal2 s 110404 -480 110516 240 8 la_data_out[1]
port 190 nsew signal output
rlabel metal2 s 164668 -480 164780 240 8 la_data_out[20]
port 191 nsew signal output
rlabel metal2 s 167524 -480 167636 240 8 la_data_out[21]
port 192 nsew signal output
rlabel metal2 s 170380 -480 170492 240 8 la_data_out[22]
port 193 nsew signal output
rlabel metal2 s 173236 -480 173348 240 8 la_data_out[23]
port 194 nsew signal output
rlabel metal2 s 176092 -480 176204 240 8 la_data_out[24]
port 195 nsew signal output
rlabel metal2 s 178948 -480 179060 240 8 la_data_out[25]
port 196 nsew signal output
rlabel metal2 s 181804 -480 181916 240 8 la_data_out[26]
port 197 nsew signal output
rlabel metal2 s 184660 -480 184772 240 8 la_data_out[27]
port 198 nsew signal output
rlabel metal2 s 187516 -480 187628 240 8 la_data_out[28]
port 199 nsew signal output
rlabel metal2 s 190372 -480 190484 240 8 la_data_out[29]
port 200 nsew signal output
rlabel metal2 s 113260 -480 113372 240 8 la_data_out[2]
port 201 nsew signal output
rlabel metal2 s 193228 -480 193340 240 8 la_data_out[30]
port 202 nsew signal output
rlabel metal2 s 196084 -480 196196 240 8 la_data_out[31]
port 203 nsew signal output
rlabel metal2 s 198940 -480 199052 240 8 la_data_out[32]
port 204 nsew signal output
rlabel metal2 s 201796 -480 201908 240 8 la_data_out[33]
port 205 nsew signal output
rlabel metal2 s 204652 -480 204764 240 8 la_data_out[34]
port 206 nsew signal output
rlabel metal2 s 207508 -480 207620 240 8 la_data_out[35]
port 207 nsew signal output
rlabel metal2 s 210364 -480 210476 240 8 la_data_out[36]
port 208 nsew signal output
rlabel metal2 s 213220 -480 213332 240 8 la_data_out[37]
port 209 nsew signal output
rlabel metal2 s 216076 -480 216188 240 8 la_data_out[38]
port 210 nsew signal output
rlabel metal2 s 218932 -480 219044 240 8 la_data_out[39]
port 211 nsew signal output
rlabel metal2 s 116116 -480 116228 240 8 la_data_out[3]
port 212 nsew signal output
rlabel metal2 s 221788 -480 221900 240 8 la_data_out[40]
port 213 nsew signal output
rlabel metal2 s 224644 -480 224756 240 8 la_data_out[41]
port 214 nsew signal output
rlabel metal2 s 227500 -480 227612 240 8 la_data_out[42]
port 215 nsew signal output
rlabel metal2 s 230356 -480 230468 240 8 la_data_out[43]
port 216 nsew signal output
rlabel metal2 s 233212 -480 233324 240 8 la_data_out[44]
port 217 nsew signal output
rlabel metal2 s 236068 -480 236180 240 8 la_data_out[45]
port 218 nsew signal output
rlabel metal2 s 238924 -480 239036 240 8 la_data_out[46]
port 219 nsew signal output
rlabel metal2 s 241780 -480 241892 240 8 la_data_out[47]
port 220 nsew signal output
rlabel metal2 s 244636 -480 244748 240 8 la_data_out[48]
port 221 nsew signal output
rlabel metal2 s 247492 -480 247604 240 8 la_data_out[49]
port 222 nsew signal output
rlabel metal2 s 118972 -480 119084 240 8 la_data_out[4]
port 223 nsew signal output
rlabel metal2 s 250348 -480 250460 240 8 la_data_out[50]
port 224 nsew signal output
rlabel metal2 s 253204 -480 253316 240 8 la_data_out[51]
port 225 nsew signal output
rlabel metal2 s 256060 -480 256172 240 8 la_data_out[52]
port 226 nsew signal output
rlabel metal2 s 258916 -480 259028 240 8 la_data_out[53]
port 227 nsew signal output
rlabel metal2 s 261772 -480 261884 240 8 la_data_out[54]
port 228 nsew signal output
rlabel metal2 s 264628 -480 264740 240 8 la_data_out[55]
port 229 nsew signal output
rlabel metal2 s 267484 -480 267596 240 8 la_data_out[56]
port 230 nsew signal output
rlabel metal2 s 270340 -480 270452 240 8 la_data_out[57]
port 231 nsew signal output
rlabel metal2 s 273196 -480 273308 240 8 la_data_out[58]
port 232 nsew signal output
rlabel metal2 s 276052 -480 276164 240 8 la_data_out[59]
port 233 nsew signal output
rlabel metal2 s 121828 -480 121940 240 8 la_data_out[5]
port 234 nsew signal output
rlabel metal2 s 278908 -480 279020 240 8 la_data_out[60]
port 235 nsew signal output
rlabel metal2 s 281764 -480 281876 240 8 la_data_out[61]
port 236 nsew signal output
rlabel metal2 s 284620 -480 284732 240 8 la_data_out[62]
port 237 nsew signal output
rlabel metal2 s 287476 -480 287588 240 8 la_data_out[63]
port 238 nsew signal output
rlabel metal2 s 124684 -480 124796 240 8 la_data_out[6]
port 239 nsew signal output
rlabel metal2 s 127540 -480 127652 240 8 la_data_out[7]
port 240 nsew signal output
rlabel metal2 s 130396 -480 130508 240 8 la_data_out[8]
port 241 nsew signal output
rlabel metal2 s 133252 -480 133364 240 8 la_data_out[9]
port 242 nsew signal output
rlabel metal2 s 108500 -480 108612 240 8 la_oenb[0]
port 243 nsew signal input
rlabel metal2 s 137060 -480 137172 240 8 la_oenb[10]
port 244 nsew signal input
rlabel metal2 s 139916 -480 140028 240 8 la_oenb[11]
port 245 nsew signal input
rlabel metal2 s 142772 -480 142884 240 8 la_oenb[12]
port 246 nsew signal input
rlabel metal2 s 145628 -480 145740 240 8 la_oenb[13]
port 247 nsew signal input
rlabel metal2 s 148484 -480 148596 240 8 la_oenb[14]
port 248 nsew signal input
rlabel metal2 s 151340 -480 151452 240 8 la_oenb[15]
port 249 nsew signal input
rlabel metal2 s 154196 -480 154308 240 8 la_oenb[16]
port 250 nsew signal input
rlabel metal2 s 157052 -480 157164 240 8 la_oenb[17]
port 251 nsew signal input
rlabel metal2 s 159908 -480 160020 240 8 la_oenb[18]
port 252 nsew signal input
rlabel metal2 s 162764 -480 162876 240 8 la_oenb[19]
port 253 nsew signal input
rlabel metal2 s 111356 -480 111468 240 8 la_oenb[1]
port 254 nsew signal input
rlabel metal2 s 165620 -480 165732 240 8 la_oenb[20]
port 255 nsew signal input
rlabel metal2 s 168476 -480 168588 240 8 la_oenb[21]
port 256 nsew signal input
rlabel metal2 s 171332 -480 171444 240 8 la_oenb[22]
port 257 nsew signal input
rlabel metal2 s 174188 -480 174300 240 8 la_oenb[23]
port 258 nsew signal input
rlabel metal2 s 177044 -480 177156 240 8 la_oenb[24]
port 259 nsew signal input
rlabel metal2 s 179900 -480 180012 240 8 la_oenb[25]
port 260 nsew signal input
rlabel metal2 s 182756 -480 182868 240 8 la_oenb[26]
port 261 nsew signal input
rlabel metal2 s 185612 -480 185724 240 8 la_oenb[27]
port 262 nsew signal input
rlabel metal2 s 188468 -480 188580 240 8 la_oenb[28]
port 263 nsew signal input
rlabel metal2 s 191324 -480 191436 240 8 la_oenb[29]
port 264 nsew signal input
rlabel metal2 s 114212 -480 114324 240 8 la_oenb[2]
port 265 nsew signal input
rlabel metal2 s 194180 -480 194292 240 8 la_oenb[30]
port 266 nsew signal input
rlabel metal2 s 197036 -480 197148 240 8 la_oenb[31]
port 267 nsew signal input
rlabel metal2 s 199892 -480 200004 240 8 la_oenb[32]
port 268 nsew signal input
rlabel metal2 s 202748 -480 202860 240 8 la_oenb[33]
port 269 nsew signal input
rlabel metal2 s 205604 -480 205716 240 8 la_oenb[34]
port 270 nsew signal input
rlabel metal2 s 208460 -480 208572 240 8 la_oenb[35]
port 271 nsew signal input
rlabel metal2 s 211316 -480 211428 240 8 la_oenb[36]
port 272 nsew signal input
rlabel metal2 s 214172 -480 214284 240 8 la_oenb[37]
port 273 nsew signal input
rlabel metal2 s 217028 -480 217140 240 8 la_oenb[38]
port 274 nsew signal input
rlabel metal2 s 219884 -480 219996 240 8 la_oenb[39]
port 275 nsew signal input
rlabel metal2 s 117068 -480 117180 240 8 la_oenb[3]
port 276 nsew signal input
rlabel metal2 s 222740 -480 222852 240 8 la_oenb[40]
port 277 nsew signal input
rlabel metal2 s 225596 -480 225708 240 8 la_oenb[41]
port 278 nsew signal input
rlabel metal2 s 228452 -480 228564 240 8 la_oenb[42]
port 279 nsew signal input
rlabel metal2 s 231308 -480 231420 240 8 la_oenb[43]
port 280 nsew signal input
rlabel metal2 s 234164 -480 234276 240 8 la_oenb[44]
port 281 nsew signal input
rlabel metal2 s 237020 -480 237132 240 8 la_oenb[45]
port 282 nsew signal input
rlabel metal2 s 239876 -480 239988 240 8 la_oenb[46]
port 283 nsew signal input
rlabel metal2 s 242732 -480 242844 240 8 la_oenb[47]
port 284 nsew signal input
rlabel metal2 s 245588 -480 245700 240 8 la_oenb[48]
port 285 nsew signal input
rlabel metal2 s 248444 -480 248556 240 8 la_oenb[49]
port 286 nsew signal input
rlabel metal2 s 119924 -480 120036 240 8 la_oenb[4]
port 287 nsew signal input
rlabel metal2 s 251300 -480 251412 240 8 la_oenb[50]
port 288 nsew signal input
rlabel metal2 s 254156 -480 254268 240 8 la_oenb[51]
port 289 nsew signal input
rlabel metal2 s 257012 -480 257124 240 8 la_oenb[52]
port 290 nsew signal input
rlabel metal2 s 259868 -480 259980 240 8 la_oenb[53]
port 291 nsew signal input
rlabel metal2 s 262724 -480 262836 240 8 la_oenb[54]
port 292 nsew signal input
rlabel metal2 s 265580 -480 265692 240 8 la_oenb[55]
port 293 nsew signal input
rlabel metal2 s 268436 -480 268548 240 8 la_oenb[56]
port 294 nsew signal input
rlabel metal2 s 271292 -480 271404 240 8 la_oenb[57]
port 295 nsew signal input
rlabel metal2 s 274148 -480 274260 240 8 la_oenb[58]
port 296 nsew signal input
rlabel metal2 s 277004 -480 277116 240 8 la_oenb[59]
port 297 nsew signal input
rlabel metal2 s 122780 -480 122892 240 8 la_oenb[5]
port 298 nsew signal input
rlabel metal2 s 279860 -480 279972 240 8 la_oenb[60]
port 299 nsew signal input
rlabel metal2 s 282716 -480 282828 240 8 la_oenb[61]
port 300 nsew signal input
rlabel metal2 s 285572 -480 285684 240 8 la_oenb[62]
port 301 nsew signal input
rlabel metal2 s 288428 -480 288540 240 8 la_oenb[63]
port 302 nsew signal input
rlabel metal2 s 125636 -480 125748 240 8 la_oenb[6]
port 303 nsew signal input
rlabel metal2 s 128492 -480 128604 240 8 la_oenb[7]
port 304 nsew signal input
rlabel metal2 s 131348 -480 131460 240 8 la_oenb[8]
port 305 nsew signal input
rlabel metal2 s 134204 -480 134316 240 8 la_oenb[9]
port 306 nsew signal input
rlabel metal2 s 289380 -480 289492 240 8 user_clock2
port 307 nsew signal input
rlabel metal2 s 290332 -480 290444 240 8 user_irq[0]
port 308 nsew signal output
rlabel metal2 s 291284 -480 291396 240 8 user_irq[1]
port 309 nsew signal output
rlabel metal2 s 292236 -480 292348 240 8 user_irq[2]
port 310 nsew signal output
rlabel metal4 s -478 -342 -168 298654 4 vdd
port 311 nsew power bidirectional
rlabel metal5 s -478 -342 298510 -32 8 vdd
port 311 nsew power bidirectional
rlabel metal5 s -478 298344 298510 298654 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 298200 -342 298510 298654 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 1577 -822 1887 299134 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 10577 -822 10887 299134 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 19577 -822 19887 299134 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 28577 -822 28887 299134 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 37577 -822 37887 299134 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 46577 -822 46887 299134 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 55577 -822 55887 299134 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 64577 -822 64887 299134 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 73577 -822 73887 299134 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 82577 -822 82887 299134 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 91577 -822 91887 299134 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 100577 -822 100887 299134 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 109577 -822 109887 299134 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 118577 -822 118887 168709 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 118577 229771 118887 299134 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 127577 -822 127887 168709 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 127577 229771 127887 299134 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 136577 -822 136887 168709 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 136577 229771 136887 299134 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 145577 -822 145887 168709 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 145577 229771 145887 299134 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 154577 -822 154887 168709 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 154577 229771 154887 299134 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 163577 -822 163887 168709 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 163577 229771 163887 299134 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 172577 -822 172887 168709 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 172577 229771 172887 299134 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 181577 -822 181887 168709 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 181577 229771 181887 299134 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 190577 -822 190887 168709 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 190577 229771 190887 299134 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 199577 -822 199887 168709 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 199577 229771 199887 299134 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 208577 -822 208887 299134 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 217577 -822 217887 299134 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 226577 -822 226887 299134 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 235577 -822 235887 299134 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 244577 -822 244887 299134 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 253577 -822 253887 299134 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 262577 -822 262887 299134 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 271577 -822 271887 299134 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 280577 -822 280887 299134 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 289577 -822 289887 299134 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -958 1913 298990 2223 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -958 10913 298990 11223 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -958 19913 298990 20223 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -958 28913 298990 29223 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -958 37913 298990 38223 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -958 46913 298990 47223 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -958 55913 298990 56223 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -958 64913 298990 65223 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -958 73913 298990 74223 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -958 82913 298990 83223 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -958 91913 298990 92223 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -958 100913 298990 101223 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -958 109913 298990 110223 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -958 118913 298990 119223 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -958 127913 298990 128223 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -958 136913 298990 137223 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -958 145913 298990 146223 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -958 154913 298990 155223 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -958 163913 298990 164223 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -958 172913 298990 173223 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -958 181913 298990 182223 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -958 190913 298990 191223 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -958 199913 298990 200223 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -958 208913 298990 209223 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -958 217913 298990 218223 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -958 226913 298990 227223 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -958 235913 298990 236223 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -958 244913 298990 245223 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -958 253913 298990 254223 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -958 262913 298990 263223 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -958 271913 298990 272223 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -958 280913 298990 281223 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -958 289913 298990 290223 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s -958 -822 -648 299134 4 vss
port 312 nsew ground bidirectional
rlabel metal5 s -958 -822 298990 -512 8 vss
port 312 nsew ground bidirectional
rlabel metal5 s -958 298824 298990 299134 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 298680 -822 298990 299134 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 3437 -822 3747 299134 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 12437 -822 12747 299134 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 21437 -822 21747 299134 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 30437 -822 30747 299134 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 39437 -822 39747 299134 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 48437 -822 48747 299134 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 57437 -822 57747 299134 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 66437 -822 66747 299134 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 75437 -822 75747 299134 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 84437 -822 84747 299134 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 93437 -822 93747 299134 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 102437 -822 102747 299134 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 111437 -822 111747 299134 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 120437 -822 120747 168709 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 120437 229771 120747 299134 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 129437 -822 129747 168709 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 129437 229771 129747 299134 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 138437 -822 138747 168709 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 138437 229771 138747 299134 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 147437 -822 147747 168709 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 147437 229771 147747 299134 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 156437 -822 156747 168709 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 156437 229771 156747 299134 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 165437 -822 165747 168709 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 165437 229771 165747 299134 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 174437 -822 174747 168709 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 174437 229771 174747 299134 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 183437 -822 183747 168709 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 183437 229771 183747 299134 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 192437 -822 192747 168709 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 192437 229771 192747 299134 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 201437 -822 201747 168709 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 201437 229771 201747 299134 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 210437 -822 210747 299134 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 219437 -822 219747 299134 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 228437 -822 228747 299134 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 237437 -822 237747 299134 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 246437 -822 246747 299134 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 255437 -822 255747 299134 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 264437 -822 264747 299134 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 273437 -822 273747 299134 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 282437 -822 282747 299134 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 291437 -822 291747 299134 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -958 4913 298990 5223 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -958 13913 298990 14223 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -958 22913 298990 23223 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -958 31913 298990 32223 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -958 40913 298990 41223 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -958 49913 298990 50223 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -958 58913 298990 59223 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -958 67913 298990 68223 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -958 76913 298990 77223 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -958 85913 298990 86223 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -958 94913 298990 95223 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -958 103913 298990 104223 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -958 112913 298990 113223 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -958 121913 298990 122223 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -958 130913 298990 131223 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -958 139913 298990 140223 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -958 148913 298990 149223 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -958 157913 298990 158223 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -958 166913 298990 167223 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -958 175913 298990 176223 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -958 184913 298990 185223 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -958 193913 298990 194223 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -958 202913 298990 203223 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -958 211913 298990 212223 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -958 220913 298990 221223 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -958 229913 298990 230223 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -958 238913 298990 239223 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -958 247913 298990 248223 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -958 256913 298990 257223 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -958 265913 298990 266223 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -958 274913 298990 275223 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -958 283913 298990 284223 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -958 292913 298990 293223 6 vss
port 312 nsew ground bidirectional
rlabel metal2 s 5684 -480 5796 240 8 wb_clk_i
port 313 nsew signal input
rlabel metal2 s 6636 -480 6748 240 8 wb_rst_i
port 314 nsew signal input
rlabel metal2 s 7588 -480 7700 240 8 wbs_ack_o
port 315 nsew signal output
rlabel metal2 s 11396 -480 11508 240 8 wbs_adr_i[0]
port 316 nsew signal input
rlabel metal2 s 43764 -480 43876 240 8 wbs_adr_i[10]
port 317 nsew signal input
rlabel metal2 s 46620 -480 46732 240 8 wbs_adr_i[11]
port 318 nsew signal input
rlabel metal2 s 49476 -480 49588 240 8 wbs_adr_i[12]
port 319 nsew signal input
rlabel metal2 s 52332 -480 52444 240 8 wbs_adr_i[13]
port 320 nsew signal input
rlabel metal2 s 55188 -480 55300 240 8 wbs_adr_i[14]
port 321 nsew signal input
rlabel metal2 s 58044 -480 58156 240 8 wbs_adr_i[15]
port 322 nsew signal input
rlabel metal2 s 60900 -480 61012 240 8 wbs_adr_i[16]
port 323 nsew signal input
rlabel metal2 s 63756 -480 63868 240 8 wbs_adr_i[17]
port 324 nsew signal input
rlabel metal2 s 66612 -480 66724 240 8 wbs_adr_i[18]
port 325 nsew signal input
rlabel metal2 s 69468 -480 69580 240 8 wbs_adr_i[19]
port 326 nsew signal input
rlabel metal2 s 15204 -480 15316 240 8 wbs_adr_i[1]
port 327 nsew signal input
rlabel metal2 s 72324 -480 72436 240 8 wbs_adr_i[20]
port 328 nsew signal input
rlabel metal2 s 75180 -480 75292 240 8 wbs_adr_i[21]
port 329 nsew signal input
rlabel metal2 s 78036 -480 78148 240 8 wbs_adr_i[22]
port 330 nsew signal input
rlabel metal2 s 80892 -480 81004 240 8 wbs_adr_i[23]
port 331 nsew signal input
rlabel metal2 s 83748 -480 83860 240 8 wbs_adr_i[24]
port 332 nsew signal input
rlabel metal2 s 86604 -480 86716 240 8 wbs_adr_i[25]
port 333 nsew signal input
rlabel metal2 s 89460 -480 89572 240 8 wbs_adr_i[26]
port 334 nsew signal input
rlabel metal2 s 92316 -480 92428 240 8 wbs_adr_i[27]
port 335 nsew signal input
rlabel metal2 s 95172 -480 95284 240 8 wbs_adr_i[28]
port 336 nsew signal input
rlabel metal2 s 98028 -480 98140 240 8 wbs_adr_i[29]
port 337 nsew signal input
rlabel metal2 s 19012 -480 19124 240 8 wbs_adr_i[2]
port 338 nsew signal input
rlabel metal2 s 100884 -480 100996 240 8 wbs_adr_i[30]
port 339 nsew signal input
rlabel metal2 s 103740 -480 103852 240 8 wbs_adr_i[31]
port 340 nsew signal input
rlabel metal2 s 22820 -480 22932 240 8 wbs_adr_i[3]
port 341 nsew signal input
rlabel metal2 s 26628 -480 26740 240 8 wbs_adr_i[4]
port 342 nsew signal input
rlabel metal2 s 29484 -480 29596 240 8 wbs_adr_i[5]
port 343 nsew signal input
rlabel metal2 s 32340 -480 32452 240 8 wbs_adr_i[6]
port 344 nsew signal input
rlabel metal2 s 35196 -480 35308 240 8 wbs_adr_i[7]
port 345 nsew signal input
rlabel metal2 s 38052 -480 38164 240 8 wbs_adr_i[8]
port 346 nsew signal input
rlabel metal2 s 40908 -480 41020 240 8 wbs_adr_i[9]
port 347 nsew signal input
rlabel metal2 s 8540 -480 8652 240 8 wbs_cyc_i
port 348 nsew signal input
rlabel metal2 s 12348 -480 12460 240 8 wbs_dat_i[0]
port 349 nsew signal input
rlabel metal2 s 44716 -480 44828 240 8 wbs_dat_i[10]
port 350 nsew signal input
rlabel metal2 s 47572 -480 47684 240 8 wbs_dat_i[11]
port 351 nsew signal input
rlabel metal2 s 50428 -480 50540 240 8 wbs_dat_i[12]
port 352 nsew signal input
rlabel metal2 s 53284 -480 53396 240 8 wbs_dat_i[13]
port 353 nsew signal input
rlabel metal2 s 56140 -480 56252 240 8 wbs_dat_i[14]
port 354 nsew signal input
rlabel metal2 s 58996 -480 59108 240 8 wbs_dat_i[15]
port 355 nsew signal input
rlabel metal2 s 61852 -480 61964 240 8 wbs_dat_i[16]
port 356 nsew signal input
rlabel metal2 s 64708 -480 64820 240 8 wbs_dat_i[17]
port 357 nsew signal input
rlabel metal2 s 67564 -480 67676 240 8 wbs_dat_i[18]
port 358 nsew signal input
rlabel metal2 s 70420 -480 70532 240 8 wbs_dat_i[19]
port 359 nsew signal input
rlabel metal2 s 16156 -480 16268 240 8 wbs_dat_i[1]
port 360 nsew signal input
rlabel metal2 s 73276 -480 73388 240 8 wbs_dat_i[20]
port 361 nsew signal input
rlabel metal2 s 76132 -480 76244 240 8 wbs_dat_i[21]
port 362 nsew signal input
rlabel metal2 s 78988 -480 79100 240 8 wbs_dat_i[22]
port 363 nsew signal input
rlabel metal2 s 81844 -480 81956 240 8 wbs_dat_i[23]
port 364 nsew signal input
rlabel metal2 s 84700 -480 84812 240 8 wbs_dat_i[24]
port 365 nsew signal input
rlabel metal2 s 87556 -480 87668 240 8 wbs_dat_i[25]
port 366 nsew signal input
rlabel metal2 s 90412 -480 90524 240 8 wbs_dat_i[26]
port 367 nsew signal input
rlabel metal2 s 93268 -480 93380 240 8 wbs_dat_i[27]
port 368 nsew signal input
rlabel metal2 s 96124 -480 96236 240 8 wbs_dat_i[28]
port 369 nsew signal input
rlabel metal2 s 98980 -480 99092 240 8 wbs_dat_i[29]
port 370 nsew signal input
rlabel metal2 s 19964 -480 20076 240 8 wbs_dat_i[2]
port 371 nsew signal input
rlabel metal2 s 101836 -480 101948 240 8 wbs_dat_i[30]
port 372 nsew signal input
rlabel metal2 s 104692 -480 104804 240 8 wbs_dat_i[31]
port 373 nsew signal input
rlabel metal2 s 23772 -480 23884 240 8 wbs_dat_i[3]
port 374 nsew signal input
rlabel metal2 s 27580 -480 27692 240 8 wbs_dat_i[4]
port 375 nsew signal input
rlabel metal2 s 30436 -480 30548 240 8 wbs_dat_i[5]
port 376 nsew signal input
rlabel metal2 s 33292 -480 33404 240 8 wbs_dat_i[6]
port 377 nsew signal input
rlabel metal2 s 36148 -480 36260 240 8 wbs_dat_i[7]
port 378 nsew signal input
rlabel metal2 s 39004 -480 39116 240 8 wbs_dat_i[8]
port 379 nsew signal input
rlabel metal2 s 41860 -480 41972 240 8 wbs_dat_i[9]
port 380 nsew signal input
rlabel metal2 s 13300 -480 13412 240 8 wbs_dat_o[0]
port 381 nsew signal output
rlabel metal2 s 45668 -480 45780 240 8 wbs_dat_o[10]
port 382 nsew signal output
rlabel metal2 s 48524 -480 48636 240 8 wbs_dat_o[11]
port 383 nsew signal output
rlabel metal2 s 51380 -480 51492 240 8 wbs_dat_o[12]
port 384 nsew signal output
rlabel metal2 s 54236 -480 54348 240 8 wbs_dat_o[13]
port 385 nsew signal output
rlabel metal2 s 57092 -480 57204 240 8 wbs_dat_o[14]
port 386 nsew signal output
rlabel metal2 s 59948 -480 60060 240 8 wbs_dat_o[15]
port 387 nsew signal output
rlabel metal2 s 62804 -480 62916 240 8 wbs_dat_o[16]
port 388 nsew signal output
rlabel metal2 s 65660 -480 65772 240 8 wbs_dat_o[17]
port 389 nsew signal output
rlabel metal2 s 68516 -480 68628 240 8 wbs_dat_o[18]
port 390 nsew signal output
rlabel metal2 s 71372 -480 71484 240 8 wbs_dat_o[19]
port 391 nsew signal output
rlabel metal2 s 17108 -480 17220 240 8 wbs_dat_o[1]
port 392 nsew signal output
rlabel metal2 s 74228 -480 74340 240 8 wbs_dat_o[20]
port 393 nsew signal output
rlabel metal2 s 77084 -480 77196 240 8 wbs_dat_o[21]
port 394 nsew signal output
rlabel metal2 s 79940 -480 80052 240 8 wbs_dat_o[22]
port 395 nsew signal output
rlabel metal2 s 82796 -480 82908 240 8 wbs_dat_o[23]
port 396 nsew signal output
rlabel metal2 s 85652 -480 85764 240 8 wbs_dat_o[24]
port 397 nsew signal output
rlabel metal2 s 88508 -480 88620 240 8 wbs_dat_o[25]
port 398 nsew signal output
rlabel metal2 s 91364 -480 91476 240 8 wbs_dat_o[26]
port 399 nsew signal output
rlabel metal2 s 94220 -480 94332 240 8 wbs_dat_o[27]
port 400 nsew signal output
rlabel metal2 s 97076 -480 97188 240 8 wbs_dat_o[28]
port 401 nsew signal output
rlabel metal2 s 99932 -480 100044 240 8 wbs_dat_o[29]
port 402 nsew signal output
rlabel metal2 s 20916 -480 21028 240 8 wbs_dat_o[2]
port 403 nsew signal output
rlabel metal2 s 102788 -480 102900 240 8 wbs_dat_o[30]
port 404 nsew signal output
rlabel metal2 s 105644 -480 105756 240 8 wbs_dat_o[31]
port 405 nsew signal output
rlabel metal2 s 24724 -480 24836 240 8 wbs_dat_o[3]
port 406 nsew signal output
rlabel metal2 s 28532 -480 28644 240 8 wbs_dat_o[4]
port 407 nsew signal output
rlabel metal2 s 31388 -480 31500 240 8 wbs_dat_o[5]
port 408 nsew signal output
rlabel metal2 s 34244 -480 34356 240 8 wbs_dat_o[6]
port 409 nsew signal output
rlabel metal2 s 37100 -480 37212 240 8 wbs_dat_o[7]
port 410 nsew signal output
rlabel metal2 s 39956 -480 40068 240 8 wbs_dat_o[8]
port 411 nsew signal output
rlabel metal2 s 42812 -480 42924 240 8 wbs_dat_o[9]
port 412 nsew signal output
rlabel metal2 s 14252 -480 14364 240 8 wbs_sel_i[0]
port 413 nsew signal input
rlabel metal2 s 18060 -480 18172 240 8 wbs_sel_i[1]
port 414 nsew signal input
rlabel metal2 s 21868 -480 21980 240 8 wbs_sel_i[2]
port 415 nsew signal input
rlabel metal2 s 25676 -480 25788 240 8 wbs_sel_i[3]
port 416 nsew signal input
rlabel metal2 s 9492 -480 9604 240 8 wbs_stb_i
port 417 nsew signal input
rlabel metal2 s 10444 -480 10556 240 8 wbs_we_i
port 418 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 298020 298020
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 16121056
string GDS_FILE /run/media/tholin/Data/Projects/MPW/AS2650/openlane/user_project_wrapper/runs/23_05_18_17_20/results/signoff/user_project_wrapper.magic.gds
string GDS_START 13493438
<< end >>

