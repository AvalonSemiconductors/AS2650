// This is the unpowered netlist.
module wrapped_as2650 (wb_clk_i,
    io_in,
    io_oeb,
    io_out);
 input wb_clk_i;
 input [37:0] io_in;
 output [37:0] io_oeb;
 output [37:0] io_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire _2933_;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire _2945_;
 wire _2946_;
 wire _2947_;
 wire _2948_;
 wire _2949_;
 wire _2950_;
 wire _2951_;
 wire _2952_;
 wire _2953_;
 wire _2954_;
 wire _2955_;
 wire _2956_;
 wire _2957_;
 wire _2958_;
 wire _2959_;
 wire _2960_;
 wire _2961_;
 wire _2962_;
 wire _2963_;
 wire _2964_;
 wire _2965_;
 wire _2966_;
 wire _2967_;
 wire _2968_;
 wire _2969_;
 wire _2970_;
 wire _2971_;
 wire _2972_;
 wire _2973_;
 wire _2974_;
 wire _2975_;
 wire _2976_;
 wire _2977_;
 wire _2978_;
 wire _2979_;
 wire _2980_;
 wire _2981_;
 wire _2982_;
 wire _2983_;
 wire _2984_;
 wire _2985_;
 wire _2986_;
 wire _2987_;
 wire _2988_;
 wire _2989_;
 wire _2990_;
 wire _2991_;
 wire _2992_;
 wire _2993_;
 wire _2994_;
 wire _2995_;
 wire _2996_;
 wire _2997_;
 wire _2998_;
 wire _2999_;
 wire _3000_;
 wire _3001_;
 wire _3002_;
 wire _3003_;
 wire _3004_;
 wire _3005_;
 wire _3006_;
 wire _3007_;
 wire _3008_;
 wire _3009_;
 wire _3010_;
 wire _3011_;
 wire _3012_;
 wire _3013_;
 wire _3014_;
 wire _3015_;
 wire _3016_;
 wire _3017_;
 wire _3018_;
 wire _3019_;
 wire _3020_;
 wire _3021_;
 wire _3022_;
 wire _3023_;
 wire _3024_;
 wire _3025_;
 wire _3026_;
 wire _3027_;
 wire _3028_;
 wire _3029_;
 wire _3030_;
 wire _3031_;
 wire _3032_;
 wire _3033_;
 wire _3034_;
 wire _3035_;
 wire _3036_;
 wire _3037_;
 wire _3038_;
 wire _3039_;
 wire _3040_;
 wire _3041_;
 wire _3042_;
 wire _3043_;
 wire _3044_;
 wire _3045_;
 wire _3046_;
 wire _3047_;
 wire _3048_;
 wire _3049_;
 wire _3050_;
 wire _3051_;
 wire _3052_;
 wire _3053_;
 wire _3054_;
 wire _3055_;
 wire _3056_;
 wire _3057_;
 wire _3058_;
 wire _3059_;
 wire _3060_;
 wire _3061_;
 wire _3062_;
 wire _3063_;
 wire _3064_;
 wire _3065_;
 wire _3066_;
 wire _3067_;
 wire _3068_;
 wire _3069_;
 wire _3070_;
 wire _3071_;
 wire _3072_;
 wire _3073_;
 wire _3074_;
 wire _3075_;
 wire _3076_;
 wire _3077_;
 wire _3078_;
 wire _3079_;
 wire _3080_;
 wire _3081_;
 wire _3082_;
 wire _3083_;
 wire _3084_;
 wire _3085_;
 wire _3086_;
 wire _3087_;
 wire _3088_;
 wire _3089_;
 wire _3090_;
 wire _3091_;
 wire _3092_;
 wire _3093_;
 wire _3094_;
 wire _3095_;
 wire _3096_;
 wire _3097_;
 wire _3098_;
 wire _3099_;
 wire _3100_;
 wire _3101_;
 wire _3102_;
 wire _3103_;
 wire _3104_;
 wire _3105_;
 wire _3106_;
 wire _3107_;
 wire _3108_;
 wire _3109_;
 wire _3110_;
 wire _3111_;
 wire _3112_;
 wire _3113_;
 wire _3114_;
 wire _3115_;
 wire _3116_;
 wire _3117_;
 wire _3118_;
 wire _3119_;
 wire _3120_;
 wire _3121_;
 wire _3122_;
 wire _3123_;
 wire _3124_;
 wire _3125_;
 wire _3126_;
 wire _3127_;
 wire _3128_;
 wire _3129_;
 wire _3130_;
 wire _3131_;
 wire _3132_;
 wire _3133_;
 wire _3134_;
 wire _3135_;
 wire _3136_;
 wire _3137_;
 wire _3138_;
 wire _3139_;
 wire _3140_;
 wire _3141_;
 wire _3142_;
 wire _3143_;
 wire _3144_;
 wire _3145_;
 wire _3146_;
 wire _3147_;
 wire _3148_;
 wire _3149_;
 wire _3150_;
 wire _3151_;
 wire _3152_;
 wire _3153_;
 wire _3154_;
 wire _3155_;
 wire _3156_;
 wire _3157_;
 wire _3158_;
 wire _3159_;
 wire _3160_;
 wire _3161_;
 wire _3162_;
 wire _3163_;
 wire _3164_;
 wire _3165_;
 wire _3166_;
 wire _3167_;
 wire _3168_;
 wire _3169_;
 wire _3170_;
 wire _3171_;
 wire _3172_;
 wire _3173_;
 wire _3174_;
 wire _3175_;
 wire _3176_;
 wire _3177_;
 wire _3178_;
 wire _3179_;
 wire _3180_;
 wire _3181_;
 wire _3182_;
 wire _3183_;
 wire _3184_;
 wire _3185_;
 wire _3186_;
 wire _3187_;
 wire _3188_;
 wire _3189_;
 wire _3190_;
 wire _3191_;
 wire _3192_;
 wire _3193_;
 wire _3194_;
 wire _3195_;
 wire _3196_;
 wire _3197_;
 wire _3198_;
 wire _3199_;
 wire _3200_;
 wire _3201_;
 wire _3202_;
 wire _3203_;
 wire _3204_;
 wire _3205_;
 wire _3206_;
 wire _3207_;
 wire _3208_;
 wire _3209_;
 wire _3210_;
 wire _3211_;
 wire _3212_;
 wire _3213_;
 wire _3214_;
 wire _3215_;
 wire _3216_;
 wire _3217_;
 wire _3218_;
 wire _3219_;
 wire _3220_;
 wire _3221_;
 wire _3222_;
 wire _3223_;
 wire _3224_;
 wire _3225_;
 wire _3226_;
 wire _3227_;
 wire _3228_;
 wire _3229_;
 wire _3230_;
 wire _3231_;
 wire _3232_;
 wire _3233_;
 wire _3234_;
 wire _3235_;
 wire _3236_;
 wire _3237_;
 wire _3238_;
 wire _3239_;
 wire _3240_;
 wire _3241_;
 wire _3242_;
 wire _3243_;
 wire _3244_;
 wire _3245_;
 wire _3246_;
 wire _3247_;
 wire _3248_;
 wire _3249_;
 wire _3250_;
 wire _3251_;
 wire _3252_;
 wire _3253_;
 wire _3254_;
 wire _3255_;
 wire _3256_;
 wire _3257_;
 wire _3258_;
 wire _3259_;
 wire _3260_;
 wire _3261_;
 wire _3262_;
 wire _3263_;
 wire _3264_;
 wire _3265_;
 wire _3266_;
 wire _3267_;
 wire _3268_;
 wire _3269_;
 wire _3270_;
 wire _3271_;
 wire _3272_;
 wire _3273_;
 wire _3274_;
 wire _3275_;
 wire _3276_;
 wire _3277_;
 wire _3278_;
 wire _3279_;
 wire _3280_;
 wire _3281_;
 wire _3282_;
 wire _3283_;
 wire _3284_;
 wire _3285_;
 wire _3286_;
 wire _3287_;
 wire _3288_;
 wire _3289_;
 wire _3290_;
 wire _3291_;
 wire _3292_;
 wire _3293_;
 wire _3294_;
 wire _3295_;
 wire _3296_;
 wire _3297_;
 wire _3298_;
 wire _3299_;
 wire _3300_;
 wire _3301_;
 wire _3302_;
 wire _3303_;
 wire _3304_;
 wire _3305_;
 wire _3306_;
 wire _3307_;
 wire _3308_;
 wire _3309_;
 wire _3310_;
 wire _3311_;
 wire _3312_;
 wire _3313_;
 wire _3314_;
 wire _3315_;
 wire _3316_;
 wire _3317_;
 wire _3318_;
 wire _3319_;
 wire _3320_;
 wire _3321_;
 wire _3322_;
 wire _3323_;
 wire _3324_;
 wire _3325_;
 wire _3326_;
 wire _3327_;
 wire _3328_;
 wire _3329_;
 wire _3330_;
 wire _3331_;
 wire _3332_;
 wire _3333_;
 wire _3334_;
 wire _3335_;
 wire _3336_;
 wire _3337_;
 wire _3338_;
 wire _3339_;
 wire _3340_;
 wire _3341_;
 wire _3342_;
 wire _3343_;
 wire _3344_;
 wire _3345_;
 wire _3346_;
 wire _3347_;
 wire _3348_;
 wire _3349_;
 wire _3350_;
 wire _3351_;
 wire _3352_;
 wire _3353_;
 wire _3354_;
 wire _3355_;
 wire _3356_;
 wire _3357_;
 wire _3358_;
 wire _3359_;
 wire _3360_;
 wire _3361_;
 wire _3362_;
 wire _3363_;
 wire _3364_;
 wire _3365_;
 wire _3366_;
 wire _3367_;
 wire _3368_;
 wire _3369_;
 wire _3370_;
 wire _3371_;
 wire _3372_;
 wire _3373_;
 wire _3374_;
 wire _3375_;
 wire _3376_;
 wire _3377_;
 wire _3378_;
 wire _3379_;
 wire _3380_;
 wire _3381_;
 wire _3382_;
 wire _3383_;
 wire _3384_;
 wire _3385_;
 wire _3386_;
 wire _3387_;
 wire _3388_;
 wire _3389_;
 wire _3390_;
 wire _3391_;
 wire _3392_;
 wire _3393_;
 wire _3394_;
 wire _3395_;
 wire _3396_;
 wire _3397_;
 wire _3398_;
 wire _3399_;
 wire _3400_;
 wire _3401_;
 wire _3402_;
 wire _3403_;
 wire _3404_;
 wire _3405_;
 wire _3406_;
 wire _3407_;
 wire _3408_;
 wire _3409_;
 wire _3410_;
 wire _3411_;
 wire _3412_;
 wire _3413_;
 wire _3414_;
 wire _3415_;
 wire _3416_;
 wire _3417_;
 wire _3418_;
 wire _3419_;
 wire _3420_;
 wire _3421_;
 wire _3422_;
 wire _3423_;
 wire _3424_;
 wire _3425_;
 wire _3426_;
 wire _3427_;
 wire _3428_;
 wire _3429_;
 wire _3430_;
 wire _3431_;
 wire _3432_;
 wire _3433_;
 wire _3434_;
 wire _3435_;
 wire _3436_;
 wire _3437_;
 wire _3438_;
 wire _3439_;
 wire _3440_;
 wire _3441_;
 wire _3442_;
 wire _3443_;
 wire _3444_;
 wire _3445_;
 wire _3446_;
 wire _3447_;
 wire _3448_;
 wire _3449_;
 wire _3450_;
 wire _3451_;
 wire _3452_;
 wire _3453_;
 wire _3454_;
 wire _3455_;
 wire _3456_;
 wire _3457_;
 wire _3458_;
 wire _3459_;
 wire _3460_;
 wire _3461_;
 wire _3462_;
 wire _3463_;
 wire _3464_;
 wire _3465_;
 wire _3466_;
 wire _3467_;
 wire _3468_;
 wire _3469_;
 wire _3470_;
 wire _3471_;
 wire _3472_;
 wire _3473_;
 wire _3474_;
 wire _3475_;
 wire _3476_;
 wire _3477_;
 wire _3478_;
 wire _3479_;
 wire _3480_;
 wire _3481_;
 wire _3482_;
 wire _3483_;
 wire _3484_;
 wire _3485_;
 wire _3486_;
 wire _3487_;
 wire _3488_;
 wire _3489_;
 wire _3490_;
 wire _3491_;
 wire _3492_;
 wire _3493_;
 wire _3494_;
 wire _3495_;
 wire _3496_;
 wire _3497_;
 wire _3498_;
 wire _3499_;
 wire _3500_;
 wire _3501_;
 wire _3502_;
 wire _3503_;
 wire _3504_;
 wire _3505_;
 wire _3506_;
 wire _3507_;
 wire _3508_;
 wire _3509_;
 wire _3510_;
 wire _3511_;
 wire _3512_;
 wire _3513_;
 wire _3514_;
 wire _3515_;
 wire _3516_;
 wire _3517_;
 wire _3518_;
 wire _3519_;
 wire _3520_;
 wire _3521_;
 wire _3522_;
 wire _3523_;
 wire _3524_;
 wire _3525_;
 wire _3526_;
 wire _3527_;
 wire _3528_;
 wire _3529_;
 wire _3530_;
 wire _3531_;
 wire _3532_;
 wire _3533_;
 wire _3534_;
 wire _3535_;
 wire _3536_;
 wire _3537_;
 wire _3538_;
 wire _3539_;
 wire _3540_;
 wire _3541_;
 wire _3542_;
 wire _3543_;
 wire _3544_;
 wire _3545_;
 wire _3546_;
 wire _3547_;
 wire _3548_;
 wire _3549_;
 wire _3550_;
 wire _3551_;
 wire _3552_;
 wire _3553_;
 wire _3554_;
 wire _3555_;
 wire _3556_;
 wire _3557_;
 wire _3558_;
 wire _3559_;
 wire _3560_;
 wire _3561_;
 wire _3562_;
 wire _3563_;
 wire _3564_;
 wire _3565_;
 wire _3566_;
 wire _3567_;
 wire _3568_;
 wire _3569_;
 wire _3570_;
 wire _3571_;
 wire _3572_;
 wire _3573_;
 wire _3574_;
 wire _3575_;
 wire _3576_;
 wire _3577_;
 wire _3578_;
 wire _3579_;
 wire _3580_;
 wire _3581_;
 wire _3582_;
 wire _3583_;
 wire _3584_;
 wire _3585_;
 wire _3586_;
 wire _3587_;
 wire _3588_;
 wire _3589_;
 wire _3590_;
 wire _3591_;
 wire _3592_;
 wire _3593_;
 wire _3594_;
 wire _3595_;
 wire _3596_;
 wire _3597_;
 wire _3598_;
 wire _3599_;
 wire _3600_;
 wire _3601_;
 wire _3602_;
 wire _3603_;
 wire _3604_;
 wire _3605_;
 wire _3606_;
 wire _3607_;
 wire _3608_;
 wire _3609_;
 wire _3610_;
 wire _3611_;
 wire _3612_;
 wire _3613_;
 wire _3614_;
 wire _3615_;
 wire _3616_;
 wire _3617_;
 wire _3618_;
 wire _3619_;
 wire _3620_;
 wire _3621_;
 wire _3622_;
 wire _3623_;
 wire _3624_;
 wire _3625_;
 wire _3626_;
 wire _3627_;
 wire _3628_;
 wire _3629_;
 wire _3630_;
 wire _3631_;
 wire _3632_;
 wire _3633_;
 wire _3634_;
 wire _3635_;
 wire _3636_;
 wire _3637_;
 wire _3638_;
 wire _3639_;
 wire _3640_;
 wire _3641_;
 wire _3642_;
 wire _3643_;
 wire _3644_;
 wire _3645_;
 wire _3646_;
 wire _3647_;
 wire _3648_;
 wire _3649_;
 wire _3650_;
 wire _3651_;
 wire _3652_;
 wire _3653_;
 wire _3654_;
 wire _3655_;
 wire _3656_;
 wire _3657_;
 wire _3658_;
 wire _3659_;
 wire _3660_;
 wire _3661_;
 wire _3662_;
 wire _3663_;
 wire _3664_;
 wire _3665_;
 wire _3666_;
 wire _3667_;
 wire _3668_;
 wire _3669_;
 wire _3670_;
 wire _3671_;
 wire _3672_;
 wire _3673_;
 wire _3674_;
 wire _3675_;
 wire _3676_;
 wire _3677_;
 wire _3678_;
 wire _3679_;
 wire _3680_;
 wire _3681_;
 wire _3682_;
 wire _3683_;
 wire _3684_;
 wire _3685_;
 wire _3686_;
 wire _3687_;
 wire _3688_;
 wire _3689_;
 wire _3690_;
 wire _3691_;
 wire _3692_;
 wire _3693_;
 wire _3694_;
 wire _3695_;
 wire _3696_;
 wire _3697_;
 wire _3698_;
 wire _3699_;
 wire _3700_;
 wire _3701_;
 wire _3702_;
 wire _3703_;
 wire _3704_;
 wire _3705_;
 wire _3706_;
 wire _3707_;
 wire _3708_;
 wire _3709_;
 wire _3710_;
 wire _3711_;
 wire _3712_;
 wire _3713_;
 wire _3714_;
 wire _3715_;
 wire _3716_;
 wire _3717_;
 wire _3718_;
 wire _3719_;
 wire _3720_;
 wire _3721_;
 wire _3722_;
 wire _3723_;
 wire _3724_;
 wire _3725_;
 wire _3726_;
 wire _3727_;
 wire _3728_;
 wire _3729_;
 wire _3730_;
 wire _3731_;
 wire _3732_;
 wire _3733_;
 wire _3734_;
 wire _3735_;
 wire _3736_;
 wire _3737_;
 wire _3738_;
 wire _3739_;
 wire _3740_;
 wire _3741_;
 wire _3742_;
 wire _3743_;
 wire _3744_;
 wire _3745_;
 wire _3746_;
 wire _3747_;
 wire _3748_;
 wire _3749_;
 wire _3750_;
 wire _3751_;
 wire _3752_;
 wire _3753_;
 wire _3754_;
 wire _3755_;
 wire _3756_;
 wire _3757_;
 wire _3758_;
 wire _3759_;
 wire _3760_;
 wire _3761_;
 wire _3762_;
 wire _3763_;
 wire _3764_;
 wire _3765_;
 wire _3766_;
 wire _3767_;
 wire _3768_;
 wire _3769_;
 wire _3770_;
 wire _3771_;
 wire _3772_;
 wire _3773_;
 wire _3774_;
 wire _3775_;
 wire _3776_;
 wire _3777_;
 wire _3778_;
 wire _3779_;
 wire _3780_;
 wire _3781_;
 wire _3782_;
 wire _3783_;
 wire _3784_;
 wire _3785_;
 wire _3786_;
 wire _3787_;
 wire _3788_;
 wire _3789_;
 wire _3790_;
 wire _3791_;
 wire _3792_;
 wire _3793_;
 wire _3794_;
 wire _3795_;
 wire _3796_;
 wire _3797_;
 wire _3798_;
 wire _3799_;
 wire _3800_;
 wire _3801_;
 wire _3802_;
 wire _3803_;
 wire _3804_;
 wire _3805_;
 wire _3806_;
 wire _3807_;
 wire _3808_;
 wire _3809_;
 wire _3810_;
 wire _3811_;
 wire _3812_;
 wire _3813_;
 wire _3814_;
 wire _3815_;
 wire _3816_;
 wire _3817_;
 wire _3818_;
 wire _3819_;
 wire _3820_;
 wire _3821_;
 wire _3822_;
 wire _3823_;
 wire _3824_;
 wire _3825_;
 wire _3826_;
 wire _3827_;
 wire _3828_;
 wire _3829_;
 wire _3830_;
 wire _3831_;
 wire _3832_;
 wire _3833_;
 wire _3834_;
 wire _3835_;
 wire _3836_;
 wire _3837_;
 wire _3838_;
 wire _3839_;
 wire _3840_;
 wire _3841_;
 wire _3842_;
 wire _3843_;
 wire _3844_;
 wire _3845_;
 wire _3846_;
 wire _3847_;
 wire _3848_;
 wire _3849_;
 wire _3850_;
 wire _3851_;
 wire _3852_;
 wire _3853_;
 wire _3854_;
 wire _3855_;
 wire _3856_;
 wire _3857_;
 wire _3858_;
 wire _3859_;
 wire _3860_;
 wire _3861_;
 wire _3862_;
 wire _3863_;
 wire _3864_;
 wire _3865_;
 wire _3866_;
 wire _3867_;
 wire _3868_;
 wire _3869_;
 wire _3870_;
 wire _3871_;
 wire _3872_;
 wire _3873_;
 wire _3874_;
 wire _3875_;
 wire _3876_;
 wire _3877_;
 wire _3878_;
 wire _3879_;
 wire _3880_;
 wire _3881_;
 wire _3882_;
 wire _3883_;
 wire _3884_;
 wire _3885_;
 wire _3886_;
 wire _3887_;
 wire _3888_;
 wire _3889_;
 wire _3890_;
 wire _3891_;
 wire _3892_;
 wire _3893_;
 wire _3894_;
 wire _3895_;
 wire _3896_;
 wire _3897_;
 wire _3898_;
 wire _3899_;
 wire _3900_;
 wire _3901_;
 wire _3902_;
 wire _3903_;
 wire _3904_;
 wire _3905_;
 wire _3906_;
 wire _3907_;
 wire _3908_;
 wire _3909_;
 wire _3910_;
 wire _3911_;
 wire _3912_;
 wire _3913_;
 wire _3914_;
 wire _3915_;
 wire _3916_;
 wire _3917_;
 wire _3918_;
 wire _3919_;
 wire _3920_;
 wire _3921_;
 wire _3922_;
 wire _3923_;
 wire _3924_;
 wire _3925_;
 wire _3926_;
 wire _3927_;
 wire _3928_;
 wire _3929_;
 wire _3930_;
 wire _3931_;
 wire _3932_;
 wire _3933_;
 wire _3934_;
 wire _3935_;
 wire _3936_;
 wire _3937_;
 wire _3938_;
 wire _3939_;
 wire _3940_;
 wire _3941_;
 wire _3942_;
 wire _3943_;
 wire _3944_;
 wire _3945_;
 wire _3946_;
 wire _3947_;
 wire _3948_;
 wire _3949_;
 wire _3950_;
 wire _3951_;
 wire _3952_;
 wire _3953_;
 wire _3954_;
 wire _3955_;
 wire _3956_;
 wire _3957_;
 wire _3958_;
 wire _3959_;
 wire _3960_;
 wire _3961_;
 wire _3962_;
 wire _3963_;
 wire _3964_;
 wire _3965_;
 wire _3966_;
 wire _3967_;
 wire _3968_;
 wire _3969_;
 wire _3970_;
 wire _3971_;
 wire _3972_;
 wire _3973_;
 wire _3974_;
 wire _3975_;
 wire _3976_;
 wire _3977_;
 wire _3978_;
 wire _3979_;
 wire _3980_;
 wire _3981_;
 wire _3982_;
 wire _3983_;
 wire _3984_;
 wire _3985_;
 wire _3986_;
 wire _3987_;
 wire _3988_;
 wire _3989_;
 wire _3990_;
 wire _3991_;
 wire _3992_;
 wire _3993_;
 wire _3994_;
 wire _3995_;
 wire _3996_;
 wire _3997_;
 wire _3998_;
 wire _3999_;
 wire _4000_;
 wire _4001_;
 wire _4002_;
 wire _4003_;
 wire _4004_;
 wire _4005_;
 wire _4006_;
 wire _4007_;
 wire _4008_;
 wire _4009_;
 wire _4010_;
 wire _4011_;
 wire _4012_;
 wire _4013_;
 wire _4014_;
 wire _4015_;
 wire _4016_;
 wire _4017_;
 wire _4018_;
 wire _4019_;
 wire _4020_;
 wire _4021_;
 wire _4022_;
 wire _4023_;
 wire _4024_;
 wire _4025_;
 wire _4026_;
 wire _4027_;
 wire _4028_;
 wire _4029_;
 wire _4030_;
 wire _4031_;
 wire _4032_;
 wire _4033_;
 wire _4034_;
 wire _4035_;
 wire _4036_;
 wire _4037_;
 wire _4038_;
 wire _4039_;
 wire _4040_;
 wire _4041_;
 wire _4042_;
 wire _4043_;
 wire _4044_;
 wire _4045_;
 wire _4046_;
 wire _4047_;
 wire _4048_;
 wire _4049_;
 wire _4050_;
 wire _4051_;
 wire _4052_;
 wire _4053_;
 wire _4054_;
 wire _4055_;
 wire _4056_;
 wire _4057_;
 wire _4058_;
 wire _4059_;
 wire _4060_;
 wire _4061_;
 wire _4062_;
 wire _4063_;
 wire _4064_;
 wire _4065_;
 wire _4066_;
 wire _4067_;
 wire _4068_;
 wire _4069_;
 wire _4070_;
 wire _4071_;
 wire _4072_;
 wire _4073_;
 wire _4074_;
 wire _4075_;
 wire _4076_;
 wire _4077_;
 wire _4078_;
 wire _4079_;
 wire _4080_;
 wire _4081_;
 wire _4082_;
 wire _4083_;
 wire _4084_;
 wire _4085_;
 wire _4086_;
 wire _4087_;
 wire _4088_;
 wire _4089_;
 wire _4090_;
 wire _4091_;
 wire _4092_;
 wire _4093_;
 wire _4094_;
 wire _4095_;
 wire _4096_;
 wire _4097_;
 wire _4098_;
 wire _4099_;
 wire _4100_;
 wire _4101_;
 wire _4102_;
 wire _4103_;
 wire _4104_;
 wire _4105_;
 wire _4106_;
 wire _4107_;
 wire _4108_;
 wire _4109_;
 wire _4110_;
 wire _4111_;
 wire _4112_;
 wire _4113_;
 wire _4114_;
 wire _4115_;
 wire _4116_;
 wire _4117_;
 wire _4118_;
 wire _4119_;
 wire _4120_;
 wire _4121_;
 wire _4122_;
 wire _4123_;
 wire _4124_;
 wire _4125_;
 wire _4126_;
 wire _4127_;
 wire _4128_;
 wire _4129_;
 wire _4130_;
 wire _4131_;
 wire _4132_;
 wire _4133_;
 wire _4134_;
 wire _4135_;
 wire _4136_;
 wire _4137_;
 wire _4138_;
 wire _4139_;
 wire _4140_;
 wire _4141_;
 wire _4142_;
 wire _4143_;
 wire _4144_;
 wire _4145_;
 wire _4146_;
 wire _4147_;
 wire _4148_;
 wire _4149_;
 wire _4150_;
 wire _4151_;
 wire _4152_;
 wire _4153_;
 wire _4154_;
 wire _4155_;
 wire _4156_;
 wire _4157_;
 wire _4158_;
 wire _4159_;
 wire _4160_;
 wire _4161_;
 wire _4162_;
 wire _4163_;
 wire _4164_;
 wire _4165_;
 wire _4166_;
 wire _4167_;
 wire _4168_;
 wire _4169_;
 wire _4170_;
 wire _4171_;
 wire _4172_;
 wire _4173_;
 wire _4174_;
 wire _4175_;
 wire _4176_;
 wire _4177_;
 wire _4178_;
 wire _4179_;
 wire _4180_;
 wire _4181_;
 wire _4182_;
 wire _4183_;
 wire _4184_;
 wire _4185_;
 wire _4186_;
 wire _4187_;
 wire _4188_;
 wire _4189_;
 wire _4190_;
 wire _4191_;
 wire _4192_;
 wire _4193_;
 wire _4194_;
 wire _4195_;
 wire _4196_;
 wire _4197_;
 wire _4198_;
 wire _4199_;
 wire _4200_;
 wire _4201_;
 wire _4202_;
 wire _4203_;
 wire _4204_;
 wire _4205_;
 wire _4206_;
 wire _4207_;
 wire _4208_;
 wire _4209_;
 wire _4210_;
 wire _4211_;
 wire _4212_;
 wire _4213_;
 wire _4214_;
 wire _4215_;
 wire _4216_;
 wire _4217_;
 wire _4218_;
 wire _4219_;
 wire _4220_;
 wire _4221_;
 wire _4222_;
 wire _4223_;
 wire _4224_;
 wire _4225_;
 wire _4226_;
 wire _4227_;
 wire _4228_;
 wire _4229_;
 wire _4230_;
 wire _4231_;
 wire _4232_;
 wire _4233_;
 wire _4234_;
 wire _4235_;
 wire _4236_;
 wire _4237_;
 wire _4238_;
 wire _4239_;
 wire _4240_;
 wire _4241_;
 wire _4242_;
 wire _4243_;
 wire _4244_;
 wire _4245_;
 wire _4246_;
 wire _4247_;
 wire _4248_;
 wire _4249_;
 wire _4250_;
 wire _4251_;
 wire _4252_;
 wire _4253_;
 wire _4254_;
 wire _4255_;
 wire _4256_;
 wire _4257_;
 wire _4258_;
 wire _4259_;
 wire _4260_;
 wire _4261_;
 wire _4262_;
 wire _4263_;
 wire _4264_;
 wire _4265_;
 wire _4266_;
 wire _4267_;
 wire _4268_;
 wire _4269_;
 wire _4270_;
 wire _4271_;
 wire _4272_;
 wire _4273_;
 wire _4274_;
 wire _4275_;
 wire _4276_;
 wire _4277_;
 wire _4278_;
 wire _4279_;
 wire _4280_;
 wire _4281_;
 wire _4282_;
 wire _4283_;
 wire _4284_;
 wire _4285_;
 wire _4286_;
 wire _4287_;
 wire _4288_;
 wire _4289_;
 wire _4290_;
 wire _4291_;
 wire _4292_;
 wire _4293_;
 wire _4294_;
 wire _4295_;
 wire _4296_;
 wire _4297_;
 wire _4298_;
 wire _4299_;
 wire _4300_;
 wire _4301_;
 wire _4302_;
 wire _4303_;
 wire _4304_;
 wire _4305_;
 wire _4306_;
 wire _4307_;
 wire _4308_;
 wire _4309_;
 wire _4310_;
 wire _4311_;
 wire _4312_;
 wire _4313_;
 wire _4314_;
 wire _4315_;
 wire _4316_;
 wire _4317_;
 wire _4318_;
 wire _4319_;
 wire _4320_;
 wire _4321_;
 wire _4322_;
 wire _4323_;
 wire _4324_;
 wire _4325_;
 wire _4326_;
 wire _4327_;
 wire _4328_;
 wire _4329_;
 wire _4330_;
 wire _4331_;
 wire _4332_;
 wire _4333_;
 wire _4334_;
 wire _4335_;
 wire _4336_;
 wire _4337_;
 wire _4338_;
 wire _4339_;
 wire _4340_;
 wire _4341_;
 wire _4342_;
 wire _4343_;
 wire _4344_;
 wire _4345_;
 wire _4346_;
 wire _4347_;
 wire _4348_;
 wire _4349_;
 wire _4350_;
 wire _4351_;
 wire _4352_;
 wire _4353_;
 wire _4354_;
 wire _4355_;
 wire _4356_;
 wire _4357_;
 wire _4358_;
 wire _4359_;
 wire _4360_;
 wire _4361_;
 wire _4362_;
 wire _4363_;
 wire _4364_;
 wire _4365_;
 wire _4366_;
 wire _4367_;
 wire _4368_;
 wire _4369_;
 wire _4370_;
 wire _4371_;
 wire _4372_;
 wire _4373_;
 wire _4374_;
 wire _4375_;
 wire _4376_;
 wire _4377_;
 wire _4378_;
 wire _4379_;
 wire _4380_;
 wire _4381_;
 wire _4382_;
 wire _4383_;
 wire _4384_;
 wire _4385_;
 wire _4386_;
 wire _4387_;
 wire _4388_;
 wire _4389_;
 wire _4390_;
 wire _4391_;
 wire _4392_;
 wire _4393_;
 wire _4394_;
 wire _4395_;
 wire _4396_;
 wire _4397_;
 wire _4398_;
 wire _4399_;
 wire _4400_;
 wire _4401_;
 wire _4402_;
 wire _4403_;
 wire _4404_;
 wire _4405_;
 wire _4406_;
 wire _4407_;
 wire _4408_;
 wire _4409_;
 wire _4410_;
 wire _4411_;
 wire _4412_;
 wire _4413_;
 wire _4414_;
 wire _4415_;
 wire _4416_;
 wire _4417_;
 wire _4418_;
 wire _4419_;
 wire _4420_;
 wire _4421_;
 wire _4422_;
 wire _4423_;
 wire _4424_;
 wire _4425_;
 wire _4426_;
 wire _4427_;
 wire _4428_;
 wire _4429_;
 wire _4430_;
 wire _4431_;
 wire _4432_;
 wire _4433_;
 wire _4434_;
 wire _4435_;
 wire _4436_;
 wire _4437_;
 wire _4438_;
 wire _4439_;
 wire _4440_;
 wire _4441_;
 wire _4442_;
 wire _4443_;
 wire _4444_;
 wire _4445_;
 wire _4446_;
 wire _4447_;
 wire _4448_;
 wire _4449_;
 wire _4450_;
 wire \as2650.addr_buff[0] ;
 wire \as2650.addr_buff[1] ;
 wire \as2650.addr_buff[2] ;
 wire \as2650.addr_buff[3] ;
 wire \as2650.addr_buff[4] ;
 wire \as2650.addr_buff[5] ;
 wire \as2650.addr_buff[6] ;
 wire \as2650.addr_buff[7] ;
 wire \as2650.alu_op[0] ;
 wire \as2650.alu_op[1] ;
 wire \as2650.alu_op[2] ;
 wire \as2650.carry ;
 wire \as2650.cycle[0] ;
 wire \as2650.cycle[10] ;
 wire \as2650.cycle[11] ;
 wire \as2650.cycle[12] ;
 wire \as2650.cycle[13] ;
 wire \as2650.cycle[1] ;
 wire \as2650.cycle[2] ;
 wire \as2650.cycle[3] ;
 wire \as2650.cycle[4] ;
 wire \as2650.cycle[5] ;
 wire \as2650.cycle[6] ;
 wire \as2650.cycle[7] ;
 wire \as2650.cycle[8] ;
 wire \as2650.cycle[9] ;
 wire \as2650.halted ;
 wire \as2650.holding_reg[0] ;
 wire \as2650.holding_reg[1] ;
 wire \as2650.holding_reg[2] ;
 wire \as2650.holding_reg[3] ;
 wire \as2650.holding_reg[4] ;
 wire \as2650.holding_reg[5] ;
 wire \as2650.holding_reg[6] ;
 wire \as2650.holding_reg[7] ;
 wire \as2650.idx_ctrl[0] ;
 wire \as2650.idx_ctrl[1] ;
 wire \as2650.ins_reg[0] ;
 wire \as2650.ins_reg[1] ;
 wire \as2650.ins_reg[2] ;
 wire \as2650.ins_reg[3] ;
 wire \as2650.ins_reg[4] ;
 wire \as2650.overflow ;
 wire \as2650.pc[0] ;
 wire \as2650.pc[10] ;
 wire \as2650.pc[11] ;
 wire \as2650.pc[12] ;
 wire \as2650.pc[13] ;
 wire \as2650.pc[14] ;
 wire \as2650.pc[1] ;
 wire \as2650.pc[2] ;
 wire \as2650.pc[3] ;
 wire \as2650.pc[4] ;
 wire \as2650.pc[5] ;
 wire \as2650.pc[6] ;
 wire \as2650.pc[7] ;
 wire \as2650.pc[8] ;
 wire \as2650.pc[9] ;
 wire \as2650.psl[1] ;
 wire \as2650.psl[3] ;
 wire \as2650.psl[4] ;
 wire \as2650.psl[5] ;
 wire \as2650.psl[6] ;
 wire \as2650.psl[7] ;
 wire \as2650.psu[0] ;
 wire \as2650.psu[1] ;
 wire \as2650.psu[2] ;
 wire \as2650.psu[3] ;
 wire \as2650.psu[4] ;
 wire \as2650.psu[5] ;
 wire \as2650.psu[7] ;
 wire \as2650.r0[0] ;
 wire \as2650.r0[1] ;
 wire \as2650.r0[2] ;
 wire \as2650.r0[3] ;
 wire \as2650.r0[4] ;
 wire \as2650.r0[5] ;
 wire \as2650.r0[6] ;
 wire \as2650.r0[7] ;
 wire \as2650.r123[0][0] ;
 wire \as2650.r123[0][1] ;
 wire \as2650.r123[0][2] ;
 wire \as2650.r123[0][3] ;
 wire \as2650.r123[0][4] ;
 wire \as2650.r123[0][5] ;
 wire \as2650.r123[0][6] ;
 wire \as2650.r123[0][7] ;
 wire \as2650.r123[1][0] ;
 wire \as2650.r123[1][1] ;
 wire \as2650.r123[1][2] ;
 wire \as2650.r123[1][3] ;
 wire \as2650.r123[1][4] ;
 wire \as2650.r123[1][5] ;
 wire \as2650.r123[1][6] ;
 wire \as2650.r123[1][7] ;
 wire \as2650.r123[2][0] ;
 wire \as2650.r123[2][1] ;
 wire \as2650.r123[2][2] ;
 wire \as2650.r123[2][3] ;
 wire \as2650.r123[2][4] ;
 wire \as2650.r123[2][5] ;
 wire \as2650.r123[2][6] ;
 wire \as2650.r123[2][7] ;
 wire \as2650.r123[3][0] ;
 wire \as2650.r123[3][1] ;
 wire \as2650.r123[3][2] ;
 wire \as2650.r123[3][3] ;
 wire \as2650.r123[3][4] ;
 wire \as2650.r123[3][5] ;
 wire \as2650.r123[3][6] ;
 wire \as2650.r123[3][7] ;
 wire \as2650.r123_2[0][0] ;
 wire \as2650.r123_2[0][1] ;
 wire \as2650.r123_2[0][2] ;
 wire \as2650.r123_2[0][3] ;
 wire \as2650.r123_2[0][4] ;
 wire \as2650.r123_2[0][5] ;
 wire \as2650.r123_2[0][6] ;
 wire \as2650.r123_2[0][7] ;
 wire \as2650.r123_2[1][0] ;
 wire \as2650.r123_2[1][1] ;
 wire \as2650.r123_2[1][2] ;
 wire \as2650.r123_2[1][3] ;
 wire \as2650.r123_2[1][4] ;
 wire \as2650.r123_2[1][5] ;
 wire \as2650.r123_2[1][6] ;
 wire \as2650.r123_2[1][7] ;
 wire \as2650.r123_2[2][0] ;
 wire \as2650.r123_2[2][1] ;
 wire \as2650.r123_2[2][2] ;
 wire \as2650.r123_2[2][3] ;
 wire \as2650.r123_2[2][4] ;
 wire \as2650.r123_2[2][5] ;
 wire \as2650.r123_2[2][6] ;
 wire \as2650.r123_2[2][7] ;
 wire \as2650.r123_2[3][0] ;
 wire \as2650.r123_2[3][1] ;
 wire \as2650.r123_2[3][2] ;
 wire \as2650.r123_2[3][3] ;
 wire \as2650.r123_2[3][4] ;
 wire \as2650.r123_2[3][5] ;
 wire \as2650.r123_2[3][6] ;
 wire \as2650.r123_2[3][7] ;
 wire \as2650.stack[0][0] ;
 wire \as2650.stack[0][10] ;
 wire \as2650.stack[0][11] ;
 wire \as2650.stack[0][12] ;
 wire \as2650.stack[0][13] ;
 wire \as2650.stack[0][14] ;
 wire \as2650.stack[0][1] ;
 wire \as2650.stack[0][2] ;
 wire \as2650.stack[0][3] ;
 wire \as2650.stack[0][4] ;
 wire \as2650.stack[0][5] ;
 wire \as2650.stack[0][6] ;
 wire \as2650.stack[0][7] ;
 wire \as2650.stack[0][8] ;
 wire \as2650.stack[0][9] ;
 wire \as2650.stack[1][0] ;
 wire \as2650.stack[1][10] ;
 wire \as2650.stack[1][11] ;
 wire \as2650.stack[1][12] ;
 wire \as2650.stack[1][13] ;
 wire \as2650.stack[1][14] ;
 wire \as2650.stack[1][1] ;
 wire \as2650.stack[1][2] ;
 wire \as2650.stack[1][3] ;
 wire \as2650.stack[1][4] ;
 wire \as2650.stack[1][5] ;
 wire \as2650.stack[1][6] ;
 wire \as2650.stack[1][7] ;
 wire \as2650.stack[1][8] ;
 wire \as2650.stack[1][9] ;
 wire \as2650.stack[2][0] ;
 wire \as2650.stack[2][10] ;
 wire \as2650.stack[2][11] ;
 wire \as2650.stack[2][12] ;
 wire \as2650.stack[2][13] ;
 wire \as2650.stack[2][14] ;
 wire \as2650.stack[2][1] ;
 wire \as2650.stack[2][2] ;
 wire \as2650.stack[2][3] ;
 wire \as2650.stack[2][4] ;
 wire \as2650.stack[2][5] ;
 wire \as2650.stack[2][6] ;
 wire \as2650.stack[2][7] ;
 wire \as2650.stack[2][8] ;
 wire \as2650.stack[2][9] ;
 wire \as2650.stack[3][0] ;
 wire \as2650.stack[3][10] ;
 wire \as2650.stack[3][11] ;
 wire \as2650.stack[3][12] ;
 wire \as2650.stack[3][13] ;
 wire \as2650.stack[3][14] ;
 wire \as2650.stack[3][1] ;
 wire \as2650.stack[3][2] ;
 wire \as2650.stack[3][3] ;
 wire \as2650.stack[3][4] ;
 wire \as2650.stack[3][5] ;
 wire \as2650.stack[3][6] ;
 wire \as2650.stack[3][7] ;
 wire \as2650.stack[3][8] ;
 wire \as2650.stack[3][9] ;
 wire \as2650.stack[4][0] ;
 wire \as2650.stack[4][10] ;
 wire \as2650.stack[4][11] ;
 wire \as2650.stack[4][12] ;
 wire \as2650.stack[4][13] ;
 wire \as2650.stack[4][14] ;
 wire \as2650.stack[4][1] ;
 wire \as2650.stack[4][2] ;
 wire \as2650.stack[4][3] ;
 wire \as2650.stack[4][4] ;
 wire \as2650.stack[4][5] ;
 wire \as2650.stack[4][6] ;
 wire \as2650.stack[4][7] ;
 wire \as2650.stack[4][8] ;
 wire \as2650.stack[4][9] ;
 wire \as2650.stack[5][0] ;
 wire \as2650.stack[5][10] ;
 wire \as2650.stack[5][11] ;
 wire \as2650.stack[5][12] ;
 wire \as2650.stack[5][13] ;
 wire \as2650.stack[5][14] ;
 wire \as2650.stack[5][1] ;
 wire \as2650.stack[5][2] ;
 wire \as2650.stack[5][3] ;
 wire \as2650.stack[5][4] ;
 wire \as2650.stack[5][5] ;
 wire \as2650.stack[5][6] ;
 wire \as2650.stack[5][7] ;
 wire \as2650.stack[5][8] ;
 wire \as2650.stack[5][9] ;
 wire \as2650.stack[6][0] ;
 wire \as2650.stack[6][10] ;
 wire \as2650.stack[6][11] ;
 wire \as2650.stack[6][12] ;
 wire \as2650.stack[6][13] ;
 wire \as2650.stack[6][14] ;
 wire \as2650.stack[6][1] ;
 wire \as2650.stack[6][2] ;
 wire \as2650.stack[6][3] ;
 wire \as2650.stack[6][4] ;
 wire \as2650.stack[6][5] ;
 wire \as2650.stack[6][6] ;
 wire \as2650.stack[6][7] ;
 wire \as2650.stack[6][8] ;
 wire \as2650.stack[6][9] ;
 wire \as2650.stack[7][0] ;
 wire \as2650.stack[7][10] ;
 wire \as2650.stack[7][11] ;
 wire \as2650.stack[7][12] ;
 wire \as2650.stack[7][13] ;
 wire \as2650.stack[7][14] ;
 wire \as2650.stack[7][1] ;
 wire \as2650.stack[7][2] ;
 wire \as2650.stack[7][3] ;
 wire \as2650.stack[7][4] ;
 wire \as2650.stack[7][5] ;
 wire \as2650.stack[7][6] ;
 wire \as2650.stack[7][7] ;
 wire \as2650.stack[7][8] ;
 wire \as2650.stack[7][9] ;
 wire net87;
 wire net92;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net88;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net89;
 wire net73;
 wire net74;
 wire net75;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire clknet_leaf_1_wb_clk_i;
 wire net90;
 wire net91;
 wire net76;
 wire net81;
 wire net77;
 wire net78;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net79;
 wire net80;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire clknet_leaf_2_wb_clk_i;
 wire clknet_leaf_3_wb_clk_i;
 wire clknet_leaf_4_wb_clk_i;
 wire clknet_leaf_5_wb_clk_i;
 wire clknet_leaf_6_wb_clk_i;
 wire clknet_leaf_7_wb_clk_i;
 wire clknet_leaf_9_wb_clk_i;
 wire clknet_leaf_13_wb_clk_i;
 wire clknet_leaf_14_wb_clk_i;
 wire clknet_leaf_15_wb_clk_i;
 wire clknet_leaf_16_wb_clk_i;
 wire clknet_leaf_17_wb_clk_i;
 wire clknet_leaf_18_wb_clk_i;
 wire clknet_leaf_19_wb_clk_i;
 wire clknet_leaf_20_wb_clk_i;
 wire clknet_leaf_21_wb_clk_i;
 wire clknet_leaf_22_wb_clk_i;
 wire clknet_leaf_23_wb_clk_i;
 wire clknet_leaf_24_wb_clk_i;
 wire clknet_leaf_25_wb_clk_i;
 wire clknet_leaf_27_wb_clk_i;
 wire clknet_leaf_29_wb_clk_i;
 wire clknet_leaf_30_wb_clk_i;
 wire clknet_leaf_31_wb_clk_i;
 wire clknet_leaf_32_wb_clk_i;
 wire clknet_leaf_33_wb_clk_i;
 wire clknet_leaf_34_wb_clk_i;
 wire clknet_leaf_35_wb_clk_i;
 wire clknet_leaf_36_wb_clk_i;
 wire clknet_leaf_37_wb_clk_i;
 wire clknet_leaf_38_wb_clk_i;
 wire clknet_leaf_40_wb_clk_i;
 wire clknet_leaf_41_wb_clk_i;
 wire clknet_leaf_43_wb_clk_i;
 wire clknet_leaf_44_wb_clk_i;
 wire clknet_leaf_45_wb_clk_i;
 wire clknet_leaf_46_wb_clk_i;
 wire clknet_leaf_47_wb_clk_i;
 wire clknet_leaf_48_wb_clk_i;
 wire clknet_leaf_49_wb_clk_i;
 wire clknet_leaf_50_wb_clk_i;
 wire clknet_leaf_51_wb_clk_i;
 wire clknet_leaf_52_wb_clk_i;
 wire clknet_leaf_53_wb_clk_i;
 wire clknet_leaf_54_wb_clk_i;
 wire clknet_leaf_55_wb_clk_i;
 wire clknet_leaf_56_wb_clk_i;
 wire clknet_leaf_57_wb_clk_i;
 wire clknet_leaf_58_wb_clk_i;
 wire clknet_leaf_59_wb_clk_i;
 wire clknet_leaf_60_wb_clk_i;
 wire clknet_leaf_61_wb_clk_i;
 wire clknet_leaf_63_wb_clk_i;
 wire clknet_leaf_66_wb_clk_i;
 wire clknet_leaf_67_wb_clk_i;
 wire clknet_leaf_68_wb_clk_i;
 wire clknet_leaf_69_wb_clk_i;
 wire clknet_leaf_70_wb_clk_i;
 wire clknet_leaf_71_wb_clk_i;
 wire clknet_leaf_73_wb_clk_i;
 wire clknet_leaf_74_wb_clk_i;
 wire clknet_leaf_75_wb_clk_i;
 wire clknet_leaf_76_wb_clk_i;
 wire clknet_leaf_77_wb_clk_i;
 wire clknet_leaf_78_wb_clk_i;
 wire clknet_leaf_79_wb_clk_i;
 wire clknet_leaf_80_wb_clk_i;
 wire clknet_leaf_81_wb_clk_i;
 wire clknet_leaf_82_wb_clk_i;
 wire clknet_0_wb_clk_i;
 wire clknet_3_0__leaf_wb_clk_i;
 wire clknet_3_1__leaf_wb_clk_i;
 wire clknet_3_2__leaf_wb_clk_i;
 wire clknet_3_3__leaf_wb_clk_i;
 wire clknet_3_4__leaf_wb_clk_i;
 wire clknet_3_5__leaf_wb_clk_i;
 wire clknet_3_6__leaf_wb_clk_i;
 wire clknet_3_7__leaf_wb_clk_i;
 wire clknet_opt_1_0_wb_clk_i;
 wire clknet_opt_2_0_wb_clk_i;
 wire clknet_opt_3_0_wb_clk_i;
 wire clknet_opt_4_0_wb_clk_i;

 gf180mcu_fd_sc_mcu7t5v0__inv_1 _4451_ (.I(\as2650.cycle[6] ),
    .ZN(_4045_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4452_ (.I(_4045_),
    .Z(_4046_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4453_ (.I(_4046_),
    .Z(_4047_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4454_ (.I(_4047_),
    .Z(_4048_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4455_ (.I(_4048_),
    .Z(_4049_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4456_ (.I(_4049_),
    .Z(_4050_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4457_ (.I(_4050_),
    .Z(_4051_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4458_ (.I(\as2650.ins_reg[4] ),
    .Z(_4052_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4459_ (.I(_4052_),
    .Z(_4053_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4460_ (.I(\as2650.alu_op[1] ),
    .Z(_4054_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4461_ (.I(_4054_),
    .Z(_4055_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4462_ (.A1(_4053_),
    .A2(_4055_),
    .ZN(_4056_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4463_ (.I(_4056_),
    .Z(_4057_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4464_ (.I(\as2650.ins_reg[0] ),
    .Z(_4058_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4465_ (.I(_4058_),
    .Z(_4059_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4466_ (.I(_4059_),
    .Z(_4060_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4467_ (.I(\as2650.psl[4] ),
    .Z(_4061_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4468_ (.I(_4061_),
    .Z(_4062_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4469_ (.I(_4062_),
    .Z(_4063_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4470_ (.I(_4063_),
    .Z(_4064_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4471_ (.I0(\as2650.r123[1][7] ),
    .I1(\as2650.r123[0][7] ),
    .I2(\as2650.r123_2[1][7] ),
    .I3(\as2650.r123_2[0][7] ),
    .S0(_4060_),
    .S1(_4064_),
    .Z(_4065_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4472_ (.I(\as2650.ins_reg[0] ),
    .Z(_4066_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _4473_ (.A1(_4066_),
    .A2(\as2650.ins_reg[1] ),
    .Z(_4067_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4474_ (.I(_4067_),
    .Z(_4068_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4475_ (.A1(_4065_),
    .A2(_4068_),
    .ZN(_4069_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4476_ (.A1(_4066_),
    .A2(\as2650.ins_reg[1] ),
    .Z(_4070_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4477_ (.I(_4070_),
    .Z(_4071_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4478_ (.I(_4071_),
    .Z(_4072_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4479_ (.I0(\as2650.r123[2][7] ),
    .I1(\as2650.r123_2[2][7] ),
    .S(_4064_),
    .Z(_4073_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4480_ (.A1(_4072_),
    .A2(_4073_),
    .ZN(_4074_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4481_ (.I(\as2650.r0[7] ),
    .Z(_4075_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4482_ (.I(_4075_),
    .Z(_4076_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4483_ (.A1(_4066_),
    .A2(\as2650.ins_reg[1] ),
    .ZN(_4077_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4484_ (.I(_4077_),
    .Z(_4078_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4485_ (.I(_4078_),
    .Z(_4079_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4486_ (.A1(_4076_),
    .A2(_4079_),
    .ZN(_4080_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _4487_ (.A1(_4069_),
    .A2(_4074_),
    .A3(_4080_),
    .ZN(_4081_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _4488_ (.I(_4063_),
    .ZN(_4082_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4489_ (.A1(_4082_),
    .A2(\as2650.r123_2[1][6] ),
    .Z(_4083_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4490_ (.I(\as2650.r123[1][6] ),
    .ZN(_4084_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4491_ (.I(\as2650.ins_reg[1] ),
    .Z(_4085_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4492_ (.I(_4085_),
    .ZN(_4086_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _4493_ (.A1(_4082_),
    .A2(_4084_),
    .B(_4086_),
    .C(_4059_),
    .ZN(_4087_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4494_ (.I(\as2650.psl[4] ),
    .Z(_4088_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4495_ (.I0(\as2650.r123[0][6] ),
    .I1(\as2650.r123_2[0][6] ),
    .S(_4088_),
    .Z(_4089_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4496_ (.I(_4089_),
    .Z(_4090_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4497_ (.I(_4090_),
    .Z(_4091_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4498_ (.I(_4091_),
    .Z(_4092_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4499_ (.I(_4059_),
    .ZN(_4093_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4500_ (.A1(_4093_),
    .A2(_4085_),
    .ZN(_4094_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _4501_ (.A1(_4083_),
    .A2(_4087_),
    .B1(_4092_),
    .B2(_4094_),
    .ZN(_4095_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4502_ (.I0(\as2650.r123[2][6] ),
    .I1(\as2650.r123_2[2][6] ),
    .S(_4063_),
    .Z(_4096_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4503_ (.A1(_4072_),
    .A2(_4096_),
    .ZN(_4097_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4504_ (.I(\as2650.r0[6] ),
    .Z(_4098_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4505_ (.I(_4098_),
    .Z(_4099_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4506_ (.I(_4099_),
    .Z(_4100_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4507_ (.A1(_4100_),
    .A2(_4079_),
    .ZN(_4101_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4508_ (.A1(_4095_),
    .A2(_4097_),
    .A3(_4101_),
    .Z(_4102_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4509_ (.I(_4102_),
    .Z(_4103_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4510_ (.I(_4103_),
    .Z(_4104_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4511_ (.I(\as2650.r0[5] ),
    .Z(_4105_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4512_ (.I(_4105_),
    .Z(_4106_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4513_ (.A1(_4106_),
    .A2(_4078_),
    .ZN(_4107_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4514_ (.I(_4061_),
    .Z(_4108_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4515_ (.I(_4108_),
    .Z(_4109_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4516_ (.I(_4109_),
    .Z(_4110_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4517_ (.I0(\as2650.r123[2][5] ),
    .I1(\as2650.r123_2[2][5] ),
    .S(_4110_),
    .Z(_4111_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4518_ (.A1(_4072_),
    .A2(_4111_),
    .ZN(_4112_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4519_ (.I0(\as2650.r123[1][5] ),
    .I1(\as2650.r123[0][5] ),
    .I2(\as2650.r123_2[1][5] ),
    .I3(\as2650.r123_2[0][5] ),
    .S0(_4059_),
    .S1(_4063_),
    .Z(_4113_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4520_ (.A1(_4068_),
    .A2(_4113_),
    .ZN(_4114_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4521_ (.A1(_4107_),
    .A2(_4112_),
    .A3(_4114_),
    .Z(_4115_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4522_ (.I(_4115_),
    .Z(_4116_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4523_ (.I(\as2650.r0[4] ),
    .Z(_4117_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4524_ (.I(_4117_),
    .Z(_4118_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4525_ (.A1(_4118_),
    .A2(_4078_),
    .ZN(_4119_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4526_ (.I0(\as2650.r123[2][4] ),
    .I1(\as2650.r123_2[2][4] ),
    .S(_4109_),
    .Z(_4120_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4527_ (.A1(_4071_),
    .A2(_4120_),
    .ZN(_4121_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4528_ (.I0(\as2650.r123[1][4] ),
    .I1(\as2650.r123[0][4] ),
    .I2(\as2650.r123_2[1][4] ),
    .I3(\as2650.r123_2[0][4] ),
    .S0(_4058_),
    .S1(_4110_),
    .Z(_4122_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4529_ (.A1(_4068_),
    .A2(_4122_),
    .ZN(_4123_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4530_ (.A1(_4119_),
    .A2(_4121_),
    .A3(_4123_),
    .Z(_4124_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4531_ (.I(_4124_),
    .Z(_4125_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4532_ (.I(_4125_),
    .Z(_4126_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4533_ (.I(\as2650.r0[3] ),
    .Z(_4127_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4534_ (.I(_4127_),
    .Z(_4128_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4535_ (.A1(_4128_),
    .A2(_4078_),
    .ZN(_4129_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4536_ (.I0(\as2650.r123[2][3] ),
    .I1(\as2650.r123_2[2][3] ),
    .S(_4110_),
    .Z(_4130_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4537_ (.I0(\as2650.r123[1][3] ),
    .I1(\as2650.r123[0][3] ),
    .I2(\as2650.r123_2[1][3] ),
    .I3(\as2650.r123_2[0][3] ),
    .S0(_4058_),
    .S1(_4110_),
    .Z(_4131_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _4538_ (.A1(_4071_),
    .A2(_4130_),
    .B1(_4131_),
    .B2(_4068_),
    .ZN(_4132_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4539_ (.A1(_4129_),
    .A2(_4132_),
    .ZN(_4133_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4540_ (.I(_4133_),
    .Z(_4134_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4541_ (.I0(\as2650.r123[2][2] ),
    .I1(\as2650.r123_2[2][2] ),
    .S(_4109_),
    .Z(_4135_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4542_ (.A1(_4071_),
    .A2(_4135_),
    .ZN(_4136_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4543_ (.I(_4136_),
    .Z(_4137_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4544_ (.I(\as2650.r0[2] ),
    .Z(_4138_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4545_ (.I(_4138_),
    .Z(_4139_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _4546_ (.I0(\as2650.r123[1][2] ),
    .I1(\as2650.r123[0][2] ),
    .I2(\as2650.r123_2[1][2] ),
    .I3(\as2650.r123_2[0][2] ),
    .S0(_4058_),
    .S1(_4109_),
    .Z(_4140_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _4547_ (.A1(_4139_),
    .A2(_4077_),
    .B1(_4140_),
    .B2(_4067_),
    .ZN(_4141_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4548_ (.I(_4141_),
    .Z(_4142_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4549_ (.A1(_4137_),
    .A2(_4142_),
    .ZN(_4143_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4550_ (.I(_4143_),
    .Z(_4144_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4551_ (.I0(\as2650.r123[1][1] ),
    .I1(\as2650.r123[0][1] ),
    .I2(\as2650.r123_2[1][1] ),
    .I3(\as2650.r123_2[0][1] ),
    .S0(_4066_),
    .S1(_4062_),
    .Z(_4145_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4552_ (.A1(_4067_),
    .A2(_4145_),
    .ZN(_4146_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4553_ (.I(_4146_),
    .Z(_4147_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4554_ (.I(_4147_),
    .Z(_4148_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4555_ (.I(\as2650.r0[1] ),
    .Z(_4149_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4556_ (.I(_4149_),
    .Z(_4150_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4557_ (.I0(\as2650.r123[2][1] ),
    .I1(\as2650.r123_2[2][1] ),
    .S(_4108_),
    .Z(_4151_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4558_ (.A1(_4150_),
    .A2(_4077_),
    .B1(_4151_),
    .B2(_4070_),
    .ZN(_4152_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4559_ (.I(_4152_),
    .Z(_4153_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4560_ (.I(_4153_),
    .Z(_4154_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4561_ (.A1(_4148_),
    .A2(_4154_),
    .ZN(_4155_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4562_ (.I(_4155_),
    .Z(_4156_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4563_ (.I(\as2650.alu_op[0] ),
    .Z(_4157_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _4564_ (.A1(_4052_),
    .A2(_4054_),
    .A3(\as2650.alu_op[2] ),
    .ZN(_4158_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4565_ (.I(\as2650.r0[0] ),
    .Z(_4159_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4566_ (.I(_4159_),
    .Z(_4160_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4567_ (.I0(\as2650.r123[2][0] ),
    .I1(\as2650.r123_2[2][0] ),
    .S(_4062_),
    .Z(_4161_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4568_ (.I0(\as2650.r123[1][0] ),
    .I1(\as2650.r123[0][0] ),
    .I2(\as2650.r123_2[1][0] ),
    .I3(\as2650.r123_2[0][0] ),
    .S0(\as2650.ins_reg[0] ),
    .S1(_4062_),
    .Z(_4162_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _4569_ (.A1(_4160_),
    .A2(_4077_),
    .B1(_4161_),
    .B2(_4070_),
    .C1(_4162_),
    .C2(_4067_),
    .ZN(_4163_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4570_ (.I(_4163_),
    .Z(_4164_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4571_ (.I(_4164_),
    .Z(_4165_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4572_ (.A1(_4157_),
    .A2(_4158_),
    .A3(_4165_),
    .ZN(_4166_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _4573_ (.A1(_4134_),
    .A2(_4144_),
    .A3(_4156_),
    .A4(_4166_),
    .ZN(_4167_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _4574_ (.A1(_4116_),
    .A2(_4126_),
    .A3(_4167_),
    .Z(_4168_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4575_ (.I(\as2650.ins_reg[4] ),
    .ZN(_4169_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _4576_ (.A1(\as2650.alu_op[0] ),
    .A2(\as2650.alu_op[1] ),
    .A3(\as2650.alu_op[2] ),
    .ZN(_4170_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4577_ (.A1(_4169_),
    .A2(_4170_),
    .ZN(_4171_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _4578_ (.A1(_4107_),
    .A2(_4112_),
    .A3(_4114_),
    .ZN(_4172_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4579_ (.I(_4172_),
    .Z(_4173_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4580_ (.A1(_4119_),
    .A2(_4121_),
    .A3(_4123_),
    .ZN(_4174_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4581_ (.I(_4174_),
    .Z(_4175_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4582_ (.I(_4163_),
    .Z(_4176_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _4583_ (.A1(_4147_),
    .A2(_4153_),
    .A3(_4176_),
    .ZN(_4177_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _4584_ (.A1(_4129_),
    .A2(_4132_),
    .A3(_4136_),
    .A4(_4141_),
    .ZN(_4178_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _4585_ (.A1(_4173_),
    .A2(_4175_),
    .A3(_4177_),
    .A4(_4178_),
    .ZN(_4179_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4586_ (.I(_4179_),
    .Z(_4180_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4587_ (.I(_4103_),
    .Z(_4181_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4588_ (.A1(_4171_),
    .A2(_4180_),
    .A3(_4181_),
    .ZN(_4182_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4589_ (.A1(_4104_),
    .A2(_4168_),
    .B(_4182_),
    .ZN(_4183_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4590_ (.A1(_4081_),
    .A2(_4183_),
    .Z(_4184_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _4591_ (.A1(_4095_),
    .A2(_4097_),
    .A3(_4101_),
    .ZN(_4185_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4592_ (.A1(_4171_),
    .A2(_4180_),
    .ZN(_4186_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4593_ (.A1(_4186_),
    .A2(_4168_),
    .ZN(_4187_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _4594_ (.A1(_4185_),
    .A2(_4187_),
    .Z(_4188_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4595_ (.I(_4126_),
    .Z(_4189_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4596_ (.A1(_4136_),
    .A2(_4141_),
    .Z(_4190_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4597_ (.I(_4190_),
    .Z(_4191_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4598_ (.I(_4191_),
    .Z(_4192_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4599_ (.I(_4176_),
    .Z(_4193_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4600_ (.A1(_4171_),
    .A2(_4193_),
    .ZN(_4194_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4601_ (.A1(_4155_),
    .A2(_4194_),
    .ZN(_4195_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4602_ (.A1(_4192_),
    .A2(_4195_),
    .ZN(_4196_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4603_ (.A1(_4134_),
    .A2(_4196_),
    .B(_4167_),
    .ZN(_4197_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4604_ (.A1(_4189_),
    .A2(_4197_),
    .Z(_4198_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _4605_ (.A1(_4129_),
    .A2(_4132_),
    .A3(_4137_),
    .A4(_4142_),
    .Z(_4199_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4606_ (.A1(_4126_),
    .A2(_4195_),
    .A3(_4199_),
    .ZN(_4200_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4607_ (.A1(_4171_),
    .A2(_4180_),
    .B1(_4200_),
    .B2(_4173_),
    .ZN(_4201_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4608_ (.I(_4173_),
    .Z(_4202_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4609_ (.A1(_4189_),
    .A2(_4167_),
    .ZN(_4203_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4610_ (.I0(_4201_),
    .I1(_4202_),
    .S(_4203_),
    .Z(_4204_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4611_ (.A1(_4129_),
    .A2(_4132_),
    .Z(_4205_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4612_ (.I(_4205_),
    .Z(_4206_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4613_ (.I(_4206_),
    .Z(_4207_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4614_ (.A1(_4146_),
    .A2(_4152_),
    .Z(_4208_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4615_ (.I(_4208_),
    .Z(_4209_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _4616_ (.A1(_4157_),
    .A2(_4158_),
    .A3(_4165_),
    .Z(_4210_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _4617_ (.A1(_4192_),
    .A2(_4209_),
    .A3(_4210_),
    .B(_4196_),
    .ZN(_4211_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4618_ (.A1(_4207_),
    .A2(_4211_),
    .Z(_4212_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4619_ (.A1(_4156_),
    .A2(_4166_),
    .B(_4195_),
    .ZN(_4213_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4620_ (.A1(_4144_),
    .A2(_4213_),
    .Z(_4214_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4621_ (.I(_4165_),
    .Z(_4215_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4622_ (.A1(_4158_),
    .A2(_4215_),
    .ZN(_4216_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4623_ (.A1(_4194_),
    .A2(_4210_),
    .ZN(_4217_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4624_ (.A1(_4209_),
    .A2(_4217_),
    .Z(_4218_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _4625_ (.A1(_4212_),
    .A2(_4214_),
    .A3(_4216_),
    .A4(_4218_),
    .Z(_4219_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _4626_ (.A1(_4198_),
    .A2(_4204_),
    .A3(_4219_),
    .ZN(_4220_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _4627_ (.A1(_4057_),
    .A2(_4184_),
    .A3(_4188_),
    .A4(_4220_),
    .ZN(_4221_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4628_ (.I(_4221_),
    .Z(_4222_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4629_ (.A1(\as2650.psl[7] ),
    .A2(_4085_),
    .Z(_4223_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4630_ (.A1(\as2650.psl[6] ),
    .A2(_4060_),
    .Z(_4224_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4631_ (.A1(_4223_),
    .A2(_4224_),
    .ZN(_4225_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4632_ (.I(_4169_),
    .Z(_4226_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4633_ (.I(_4054_),
    .ZN(_4227_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4634_ (.I(\as2650.alu_op[2] ),
    .Z(_4228_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4635_ (.A1(_4227_),
    .A2(_4228_),
    .ZN(_4229_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4636_ (.I(_4229_),
    .Z(_4230_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4637_ (.A1(_4226_),
    .A2(_4230_),
    .ZN(_4231_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4638_ (.I(_4072_),
    .Z(_4232_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4639_ (.A1(_4054_),
    .A2(_4228_),
    .ZN(_4233_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4640_ (.A1(_4053_),
    .A2(_4233_),
    .ZN(_4234_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4641_ (.A1(_4232_),
    .A2(_4225_),
    .A3(_4234_),
    .ZN(_4235_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _4642_ (.A1(_4225_),
    .A2(_4231_),
    .B(_4235_),
    .ZN(_4236_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _4643_ (.I(_4236_),
    .ZN(_4237_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4644_ (.I(\as2650.ins_reg[3] ),
    .Z(_4238_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4645_ (.I(_4052_),
    .Z(_4239_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4646_ (.A1(_4238_),
    .A2(_4239_),
    .ZN(_4240_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4647_ (.I(_4240_),
    .Z(_4241_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4648_ (.I(_4241_),
    .Z(_4242_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4649_ (.I(\as2650.halted ),
    .ZN(_4243_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4650_ (.I(net5),
    .ZN(_4244_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4651_ (.A1(_4243_),
    .A2(_4244_),
    .ZN(_4245_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4652_ (.I(_4245_),
    .Z(_4246_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4653_ (.A1(_4242_),
    .A2(_4246_),
    .ZN(_4247_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4654_ (.I(_4232_),
    .Z(_4248_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4655_ (.I(_4228_),
    .ZN(_4249_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4656_ (.A1(_4055_),
    .A2(_4249_),
    .ZN(_4250_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4657_ (.I(_4250_),
    .Z(_4251_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4658_ (.I(\as2650.ins_reg[3] ),
    .ZN(_4252_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4659_ (.I(_4252_),
    .Z(_4253_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4660_ (.A1(_4253_),
    .A2(_4226_),
    .ZN(_4254_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _4661_ (.A1(_4248_),
    .A2(_4251_),
    .A3(_4254_),
    .ZN(_4255_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4662_ (.I(_4255_),
    .Z(_4256_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4663_ (.A1(_4247_),
    .A2(_4256_),
    .ZN(_4257_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _4664_ (.A1(_4051_),
    .A2(_4222_),
    .A3(_4237_),
    .A4(_4257_),
    .Z(_4258_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4665_ (.I(net5),
    .Z(_4259_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4666_ (.A1(net6),
    .A2(\as2650.cycle[13] ),
    .ZN(_4260_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4667_ (.I(_4260_),
    .Z(_4261_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4668_ (.I(_4261_),
    .Z(_4262_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4669_ (.I(net6),
    .Z(_4263_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4670_ (.I(_4263_),
    .Z(_4264_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4671_ (.I(_4264_),
    .Z(_4265_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4672_ (.A1(_4265_),
    .A2(\as2650.cycle[7] ),
    .ZN(_4266_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4673_ (.I(_4266_),
    .ZN(_4267_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4674_ (.I(\as2650.ins_reg[2] ),
    .Z(_4268_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _4675_ (.I(_4268_),
    .ZN(_4269_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4676_ (.A1(_4269_),
    .A2(_4255_),
    .ZN(_4270_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4677_ (.I(_4264_),
    .Z(_4271_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4678_ (.A1(_4271_),
    .A2(\as2650.cycle[12] ),
    .ZN(_4272_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4679_ (.I(_4263_),
    .Z(_4273_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4680_ (.A1(_4273_),
    .A2(\as2650.cycle[5] ),
    .ZN(_4274_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _4681_ (.A1(_4270_),
    .A2(_4272_),
    .A3(_4274_),
    .ZN(_4275_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4682_ (.I(_4254_),
    .Z(_4276_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4683_ (.I(_4268_),
    .Z(_4277_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4684_ (.A1(_4232_),
    .A2(_4250_),
    .ZN(_4278_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4685_ (.A1(_4278_),
    .A2(_4240_),
    .ZN(_4279_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4686_ (.A1(_4277_),
    .A2(_4279_),
    .ZN(_4280_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4687_ (.A1(_4264_),
    .A2(\as2650.cycle[11] ),
    .ZN(_4281_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4688_ (.I(\as2650.cycle[5] ),
    .ZN(_4282_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _4689_ (.I(\as2650.cycle[4] ),
    .ZN(_4283_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4690_ (.A1(_4282_),
    .A2(_4283_),
    .ZN(_4284_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4691_ (.A1(_4273_),
    .A2(_4284_),
    .ZN(_4285_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _4692_ (.A1(_4276_),
    .A2(_4280_),
    .A3(_4281_),
    .A4(_4285_),
    .ZN(_4286_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4693_ (.A1(_4277_),
    .A2(_4240_),
    .ZN(_4287_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4694_ (.A1(_4232_),
    .A2(_4250_),
    .A3(_4287_),
    .ZN(_4288_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4695_ (.A1(_4267_),
    .A2(_4275_),
    .B(_4286_),
    .C(_4288_),
    .ZN(_4289_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4696_ (.I(\as2650.halted ),
    .Z(_4290_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4697_ (.A1(_4262_),
    .A2(_4289_),
    .B(_4290_),
    .ZN(_4291_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4698_ (.A1(_4259_),
    .A2(_4291_),
    .Z(_4292_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4699_ (.I(_4238_),
    .Z(_4293_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4700_ (.I(_4293_),
    .Z(_4294_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4701_ (.I(_4277_),
    .Z(_4295_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4702_ (.I(_4295_),
    .Z(_4296_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4703_ (.I(_4053_),
    .Z(_4297_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4704_ (.I(_4297_),
    .Z(_4298_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4705_ (.I(_4233_),
    .Z(_4299_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4706_ (.A1(_4296_),
    .A2(_4298_),
    .A3(_4299_),
    .ZN(_4300_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4707_ (.A1(_4294_),
    .A2(_4300_),
    .ZN(_4301_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4708_ (.I(\as2650.alu_op[0] ),
    .Z(_4302_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4709_ (.I(_4227_),
    .Z(_4303_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4710_ (.A1(_4302_),
    .A2(_4303_),
    .ZN(_4304_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4711_ (.A1(_4269_),
    .A2(_4053_),
    .A3(_4304_),
    .ZN(_4305_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4712_ (.I(_4305_),
    .Z(_4306_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4713_ (.A1(_4293_),
    .A2(_4306_),
    .ZN(_4307_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4714_ (.I(_4307_),
    .Z(_4308_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4715_ (.A1(\as2650.halted ),
    .A2(net5),
    .ZN(_4309_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4716_ (.I(_4309_),
    .Z(_4310_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4717_ (.I(_4310_),
    .Z(_4311_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4718_ (.A1(_4301_),
    .A2(_4308_),
    .B(_4311_),
    .ZN(_4312_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4719_ (.I(_4261_),
    .Z(_4313_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4720_ (.I(_4313_),
    .Z(_4314_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4721_ (.A1(_4252_),
    .A2(_4239_),
    .ZN(_4315_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4722_ (.A1(_4052_),
    .A2(_4157_),
    .ZN(_4316_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4723_ (.A1(_4268_),
    .A2(_4316_),
    .ZN(_4317_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4724_ (.A1(_4249_),
    .A2(_4317_),
    .ZN(_4318_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4725_ (.A1(_4315_),
    .A2(_4318_),
    .ZN(_4319_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4726_ (.I(_4319_),
    .Z(_4320_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4727_ (.A1(_4311_),
    .A2(_4314_),
    .A3(_4320_),
    .ZN(_4321_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4728_ (.A1(_4238_),
    .A2(_4169_),
    .ZN(_4322_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4729_ (.I(_4322_),
    .Z(_4323_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4730_ (.I(_4269_),
    .Z(_4324_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4731_ (.A1(_4324_),
    .A2(_4234_),
    .ZN(_4325_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _4732_ (.A1(_4269_),
    .A2(_4239_),
    .A3(_4157_),
    .ZN(_4326_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4733_ (.A1(_4306_),
    .A2(_4326_),
    .ZN(_4327_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4734_ (.A1(_4325_),
    .A2(_4327_),
    .ZN(_4328_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4735_ (.I(_4328_),
    .Z(_4329_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _4736_ (.A1(_4311_),
    .A2(_4262_),
    .A3(_4323_),
    .A4(_4329_),
    .ZN(_4330_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _4737_ (.A1(_4292_),
    .A2(_4312_),
    .A3(_4321_),
    .A4(_4330_),
    .ZN(_4331_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4738_ (.A1(_4264_),
    .A2(\as2650.cycle[3] ),
    .Z(_4332_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4739_ (.A1(_4263_),
    .A2(\as2650.cycle[1] ),
    .Z(_4333_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4740_ (.A1(_4332_),
    .A2(_4333_),
    .ZN(_4334_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4741_ (.I(_4334_),
    .Z(_4335_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4742_ (.I(_4335_),
    .Z(_4336_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4743_ (.I(\as2650.cycle[10] ),
    .Z(_4337_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4744_ (.A1(\as2650.cycle[2] ),
    .A2(_4337_),
    .B(_4271_),
    .ZN(_4338_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4745_ (.I(_4338_),
    .Z(_4339_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4746_ (.A1(_4336_),
    .A2(_4339_),
    .ZN(_4340_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4747_ (.I(_4226_),
    .Z(_4341_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4748_ (.I(_4341_),
    .Z(_4342_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4749_ (.I(_4244_),
    .Z(_4343_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4750_ (.A1(net6),
    .A2(\as2650.cycle[13] ),
    .Z(_4344_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4751_ (.I(_4344_),
    .Z(_4345_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4752_ (.I(_4345_),
    .Z(_4346_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4753_ (.A1(_4263_),
    .A2(\as2650.cycle[11] ),
    .Z(_4347_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4754_ (.I(_4347_),
    .Z(_4348_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4755_ (.I(_4348_),
    .Z(_4349_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4756_ (.A1(_4290_),
    .A2(_4346_),
    .A3(_4349_),
    .ZN(_4350_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _4757_ (.A1(_4342_),
    .A2(_4343_),
    .A3(_4350_),
    .ZN(_4351_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4758_ (.A1(_4340_),
    .A2(_4351_),
    .ZN(_4352_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4759_ (.I(\as2650.cycle[13] ),
    .Z(_4353_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4760_ (.I(_4353_),
    .Z(_4354_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4761_ (.A1(_4331_),
    .A2(_4352_),
    .B(_4354_),
    .ZN(_4355_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4762_ (.I(\as2650.cycle[6] ),
    .Z(_4356_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4763_ (.I(_4356_),
    .Z(_4357_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4764_ (.I(_4357_),
    .Z(_4358_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4765_ (.I(_4358_),
    .Z(_4359_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4766_ (.I(_4359_),
    .Z(_4360_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4767_ (.I(_4360_),
    .Z(_4361_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4768_ (.I(_4361_),
    .Z(_4362_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4769_ (.I(_4362_),
    .Z(_4363_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4770_ (.I(_4311_),
    .Z(_4364_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4771_ (.I(_4364_),
    .Z(_4365_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4772_ (.I(_4365_),
    .Z(_4366_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4773_ (.I(_4294_),
    .Z(_4367_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4774_ (.I(_4367_),
    .Z(_4368_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4775_ (.A1(_4293_),
    .A2(_4324_),
    .ZN(_4369_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4776_ (.I(_4369_),
    .Z(_4370_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4777_ (.I(_4315_),
    .Z(_4371_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4778_ (.I(_4093_),
    .Z(_4372_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4779_ (.A1(_4372_),
    .A2(_4086_),
    .ZN(_4373_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4780_ (.I(_4373_),
    .Z(_4374_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4781_ (.A1(\as2650.ins_reg[3] ),
    .A2(\as2650.ins_reg[2] ),
    .Z(_4375_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4782_ (.I(_4375_),
    .Z(_4376_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4783_ (.I(_4376_),
    .Z(_4377_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4784_ (.I(_4377_),
    .Z(_4378_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4785_ (.I(_4378_),
    .Z(_4379_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4786_ (.A1(_4374_),
    .A2(_4379_),
    .ZN(_4380_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4787_ (.I(_4302_),
    .Z(_4381_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4788_ (.A1(_4381_),
    .A2(_4229_),
    .ZN(_4382_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4789_ (.I(_4382_),
    .Z(_4383_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _4790_ (.A1(_4298_),
    .A2(_4380_),
    .A3(_4383_),
    .ZN(_4384_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4791_ (.A1(_4328_),
    .A2(_4384_),
    .ZN(_4385_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4792_ (.I(_4239_),
    .Z(_4386_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4793_ (.I(_4386_),
    .Z(_4387_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4794_ (.I(_4387_),
    .Z(_4388_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4795_ (.I(_4302_),
    .Z(_4389_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4796_ (.I(_4389_),
    .Z(_4390_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4797_ (.I(_4390_),
    .Z(_4391_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4798_ (.I(_4303_),
    .Z(_4392_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4799_ (.I(_4079_),
    .Z(_4393_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4800_ (.A1(\as2650.ins_reg[3] ),
    .A2(\as2650.ins_reg[2] ),
    .ZN(_4394_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4801_ (.I(_4394_),
    .Z(_4395_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4802_ (.I(_4395_),
    .Z(_4396_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4803_ (.I(_4396_),
    .Z(_4397_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4804_ (.A1(_4393_),
    .A2(_4397_),
    .ZN(_4398_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _4805_ (.A1(_4388_),
    .A2(_4391_),
    .A3(_4392_),
    .A4(_4398_),
    .ZN(_4399_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4806_ (.I(_4388_),
    .Z(_4400_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4807_ (.I(_4400_),
    .Z(_4401_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4808_ (.I(_4401_),
    .Z(_4402_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4809_ (.A1(_4371_),
    .A2(_4385_),
    .B1(_4399_),
    .B2(_4402_),
    .ZN(_4403_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4810_ (.A1(_4370_),
    .A2(_4403_),
    .ZN(_4404_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4811_ (.A1(_4295_),
    .A2(_4255_),
    .ZN(_4405_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _4812_ (.I(_4405_),
    .ZN(_4406_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4813_ (.A1(_4368_),
    .A2(_4326_),
    .B(_4404_),
    .C(_4406_),
    .ZN(_4407_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4814_ (.A1(_4363_),
    .A2(_4366_),
    .A3(_4407_),
    .ZN(_4408_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4815_ (.I(_4333_),
    .Z(_4409_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4816_ (.I(_4409_),
    .Z(_4410_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4817_ (.I(\as2650.addr_buff[7] ),
    .Z(_4411_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4818_ (.A1(_4271_),
    .A2(\as2650.cycle[10] ),
    .ZN(_4412_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4819_ (.A1(\as2650.cycle[3] ),
    .A2(_4411_),
    .A3(_4412_),
    .ZN(_4413_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4820_ (.I(net3),
    .Z(_4414_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4821_ (.I(_4414_),
    .Z(_4415_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4822_ (.A1(_4415_),
    .A2(_4409_),
    .ZN(_4416_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4823_ (.A1(_4410_),
    .A2(_4413_),
    .B(_4416_),
    .ZN(_4417_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4824_ (.A1(\as2650.cycle[9] ),
    .A2(_4335_),
    .A3(_4338_),
    .ZN(_4418_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4825_ (.I(_4249_),
    .Z(_4419_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4826_ (.A1(_4381_),
    .A2(_4303_),
    .A3(_4419_),
    .ZN(_4420_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4827_ (.A1(_4417_),
    .A2(_4418_),
    .B(_4420_),
    .C(_4351_),
    .ZN(_4421_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4828_ (.I(_4421_),
    .ZN(_4422_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4829_ (.I(_4270_),
    .Z(_4423_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4830_ (.I(_4423_),
    .Z(_4424_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4831_ (.I(_4424_),
    .Z(_4425_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4832_ (.A1(_4363_),
    .A2(_4366_),
    .A3(_4425_),
    .ZN(_4426_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _4833_ (.A1(_4355_),
    .A2(_4408_),
    .A3(_4422_),
    .A4(_4426_),
    .Z(_4427_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4834_ (.A1(_4258_),
    .A2(_4427_),
    .ZN(_0004_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4835_ (.I(_4314_),
    .Z(_4428_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4836_ (.A1(_4424_),
    .A2(_4428_),
    .ZN(_4429_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4837_ (.I(_4411_),
    .Z(_4430_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4838_ (.I(_4430_),
    .Z(_4431_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4839_ (.I(_4431_),
    .Z(_4432_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4840_ (.I(\as2650.cycle[5] ),
    .Z(_4433_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4841_ (.A1(_4265_),
    .A2(_4433_),
    .Z(_4434_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4842_ (.I(_4434_),
    .Z(_4435_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4843_ (.I(_4435_),
    .Z(_4436_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4844_ (.I(_4436_),
    .Z(_4437_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4845_ (.I(_4253_),
    .Z(_4438_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4846_ (.I(_4438_),
    .Z(_4439_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4847_ (.I(_4439_),
    .Z(_4440_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4848_ (.A1(_4296_),
    .A2(_4278_),
    .A3(_4240_),
    .ZN(_4441_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4849_ (.I(_4441_),
    .Z(_4442_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4850_ (.A1(_4440_),
    .A2(_4442_),
    .ZN(_4443_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _4851_ (.A1(_4432_),
    .A2(_4365_),
    .A3(_4437_),
    .A4(_4443_),
    .ZN(_4444_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4852_ (.I(_4323_),
    .Z(_4445_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4853_ (.A1(_4364_),
    .A2(_4445_),
    .ZN(_4446_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4854_ (.I(_4274_),
    .Z(_4447_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4855_ (.I(_4447_),
    .Z(_4448_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4856_ (.I(_4419_),
    .Z(_4449_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4857_ (.I(_4449_),
    .Z(_4450_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4858_ (.A1(_4450_),
    .A2(_4326_),
    .ZN(_0290_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4859_ (.A1(_4448_),
    .A2(_0290_),
    .ZN(_0291_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4860_ (.I(_4331_),
    .ZN(_0292_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4861_ (.A1(_4446_),
    .A2(_0291_),
    .B(_0292_),
    .ZN(_0293_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4862_ (.A1(_4352_),
    .A2(_0293_),
    .ZN(_0294_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4863_ (.I(_0294_),
    .ZN(_0295_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4864_ (.I(_0295_),
    .Z(_0296_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4865_ (.A1(\as2650.cycle[12] ),
    .A2(_0296_),
    .ZN(_0297_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4866_ (.A1(_4429_),
    .A2(_4444_),
    .B(_0297_),
    .ZN(_0003_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4867_ (.I(_4365_),
    .Z(_0298_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4868_ (.I(_4428_),
    .Z(_0299_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4869_ (.I(_0299_),
    .Z(_0300_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4870_ (.A1(_4226_),
    .A2(_4420_),
    .Z(_0301_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4871_ (.I(_0301_),
    .Z(_0302_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4872_ (.I(_0302_),
    .Z(_0303_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4873_ (.A1(_4370_),
    .A2(_0303_),
    .ZN(_0304_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4874_ (.I(_4401_),
    .Z(_0305_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4875_ (.I(_0305_),
    .Z(_0306_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4876_ (.A1(_4283_),
    .A2(_0306_),
    .ZN(_0307_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _4877_ (.A1(_0298_),
    .A2(_0300_),
    .A3(_0304_),
    .A4(_0307_),
    .ZN(_0308_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4878_ (.I(_4271_),
    .Z(_0309_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4879_ (.A1(_4433_),
    .A2(_4283_),
    .ZN(_0310_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _4880_ (.A1(_0309_),
    .A2(_4255_),
    .A3(_4313_),
    .A4(_0310_),
    .Z(_0311_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4881_ (.A1(\as2650.cycle[11] ),
    .A2(_0295_),
    .B1(_0311_),
    .B2(_4247_),
    .ZN(_0312_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4882_ (.A1(_0308_),
    .A2(_0312_),
    .ZN(_0002_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4883_ (.I(\as2650.cycle[1] ),
    .ZN(_0313_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4884_ (.I(_4332_),
    .Z(_0314_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4885_ (.A1(_0313_),
    .A2(_0314_),
    .ZN(_0315_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4886_ (.A1(_4337_),
    .A2(_0296_),
    .ZN(_0316_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4887_ (.A1(_4351_),
    .A2(_0315_),
    .B(_0316_),
    .ZN(_0001_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4888_ (.I(\as2650.cycle[9] ),
    .Z(_0317_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4889_ (.I(_0317_),
    .Z(_0318_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4890_ (.A1(_0318_),
    .A2(_0293_),
    .ZN(_0319_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4891_ (.I(_4342_),
    .Z(_0320_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4892_ (.I(_0320_),
    .Z(_0321_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4893_ (.I(_4259_),
    .Z(_0322_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4894_ (.A1(_4273_),
    .A2(\as2650.cycle[3] ),
    .ZN(_0323_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4895_ (.I(_0323_),
    .Z(_0324_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4896_ (.I(_4412_),
    .Z(_0325_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4897_ (.I(_0325_),
    .Z(_0326_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4898_ (.A1(_0324_),
    .A2(_0326_),
    .ZN(_0327_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4899_ (.A1(_0322_),
    .A2(_0327_),
    .ZN(_0328_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4900_ (.A1(\as2650.cycle[2] ),
    .A2(_4265_),
    .ZN(_0329_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4901_ (.I(_0329_),
    .Z(_0330_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4902_ (.A1(\as2650.cycle[1] ),
    .A2(_0330_),
    .ZN(_0331_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _4903_ (.A1(_0321_),
    .A2(_4350_),
    .A3(_0328_),
    .A4(_0331_),
    .ZN(_0332_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4904_ (.A1(_0319_),
    .A2(_0332_),
    .ZN(_0013_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4905_ (.I(_0322_),
    .Z(_0333_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4906_ (.I(_0333_),
    .Z(_0334_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4907_ (.I(_0334_),
    .Z(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4908_ (.I(_4243_),
    .Z(_0336_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4909_ (.I(\as2650.cycle[0] ),
    .Z(_0337_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4910_ (.I(_0337_),
    .Z(_0338_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4911_ (.I(_0338_),
    .Z(_0339_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4912_ (.I(_0339_),
    .Z(_0340_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4913_ (.I(\as2650.cycle[8] ),
    .Z(_0341_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4914_ (.I(_0341_),
    .Z(_0342_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4915_ (.A1(_0336_),
    .A2(_0309_),
    .ZN(_0343_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4916_ (.A1(_0336_),
    .A2(_0340_),
    .B1(_0342_),
    .B2(_0343_),
    .ZN(_0344_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4917_ (.A1(_0335_),
    .A2(_0344_),
    .ZN(_0012_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _4918_ (.A1(_0309_),
    .A2(_4282_),
    .A3(\as2650.cycle[12] ),
    .A4(_4270_),
    .ZN(_0345_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4919_ (.I(\as2650.cycle[7] ),
    .ZN(_0346_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _4920_ (.A1(_4354_),
    .A2(_4246_),
    .A3(_0345_),
    .B1(_0294_),
    .B2(_0346_),
    .ZN(_0011_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4921_ (.I(\as2650.cycle[8] ),
    .ZN(_0347_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4922_ (.I(_0347_),
    .Z(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4923_ (.I(_0333_),
    .Z(_0349_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4924_ (.I(_4343_),
    .Z(_0350_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4925_ (.I(_0350_),
    .Z(_0351_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4926_ (.A1(_4363_),
    .A2(_0351_),
    .ZN(_0352_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _4927_ (.A1(_0348_),
    .A2(_0349_),
    .A3(_0343_),
    .B1(_0352_),
    .B2(_0336_),
    .ZN(_0010_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4928_ (.I(_4433_),
    .Z(_0353_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4929_ (.I(_0353_),
    .Z(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4930_ (.I(_0354_),
    .Z(_0355_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4931_ (.A1(_0355_),
    .A2(_0293_),
    .ZN(_0356_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4932_ (.I(_4346_),
    .Z(_0357_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4933_ (.I(_0357_),
    .Z(_0358_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4934_ (.I(_4280_),
    .Z(_0359_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4935_ (.I(_0359_),
    .Z(_0360_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4936_ (.A1(_4400_),
    .A2(_0360_),
    .ZN(_0361_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4937_ (.A1(_0298_),
    .A2(_0358_),
    .A3(_0361_),
    .ZN(_0362_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4938_ (.A1(_4341_),
    .A2(_4304_),
    .A3(_4380_),
    .ZN(_0363_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4939_ (.A1(_4047_),
    .A2(_4388_),
    .ZN(_0364_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4940_ (.I(_0364_),
    .Z(_0365_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4941_ (.A1(_4365_),
    .A2(_0363_),
    .A3(_0365_),
    .ZN(_0366_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4942_ (.I(_4397_),
    .Z(_0367_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4943_ (.I(_0367_),
    .Z(_0368_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4944_ (.I(_0368_),
    .Z(_0369_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4945_ (.I(_4228_),
    .Z(_0370_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4946_ (.A1(_4302_),
    .A2(_4055_),
    .A3(_0370_),
    .ZN(_0371_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4947_ (.A1(_4342_),
    .A2(_0371_),
    .ZN(_0372_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4948_ (.I(_0372_),
    .Z(_0373_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4949_ (.A1(_0369_),
    .A2(_0373_),
    .ZN(_0374_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4950_ (.A1(_4296_),
    .A2(_4345_),
    .ZN(_0375_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4951_ (.I(_0375_),
    .Z(_0376_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4952_ (.I(_0376_),
    .Z(_0377_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _4953_ (.A1(_4420_),
    .A2(_0366_),
    .A3(_0374_),
    .B1(_0377_),
    .B2(_4257_),
    .ZN(_0378_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4954_ (.I(_0378_),
    .ZN(_0379_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4955_ (.I(_4445_),
    .Z(_0380_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4956_ (.I(_0290_),
    .Z(_0381_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _4957_ (.A1(_4354_),
    .A2(_0298_),
    .A3(_0380_),
    .A4(_0381_),
    .ZN(_0382_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _4958_ (.A1(_0356_),
    .A2(_0362_),
    .A3(_0379_),
    .A4(_0382_),
    .ZN(_0009_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4959_ (.I(\as2650.cycle[4] ),
    .Z(_0383_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4960_ (.A1(_0383_),
    .A2(_0293_),
    .ZN(_0384_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4961_ (.I(_4400_),
    .Z(_0385_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4962_ (.I(_0385_),
    .Z(_0386_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4963_ (.I(_0386_),
    .Z(_0387_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4964_ (.I(_0359_),
    .Z(_0388_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4965_ (.A1(_0388_),
    .A2(_4314_),
    .ZN(_0389_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4966_ (.I(net3),
    .Z(_0390_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4967_ (.I(_0390_),
    .Z(_0391_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4968_ (.I(_0391_),
    .Z(_0392_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4969_ (.I(_0392_),
    .Z(_0393_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4970_ (.I(_0393_),
    .Z(_0394_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4971_ (.I(_4443_),
    .Z(_0395_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4972_ (.A1(_4295_),
    .A2(_4261_),
    .ZN(_0396_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4973_ (.I(_0396_),
    .Z(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4974_ (.I(_0397_),
    .Z(_0398_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4975_ (.I(_0398_),
    .Z(_0399_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _4976_ (.A1(_0394_),
    .A2(_4366_),
    .A3(_0395_),
    .A4(_0399_),
    .ZN(_0400_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4977_ (.A1(_4444_),
    .A2(_0389_),
    .B(_0400_),
    .ZN(_0401_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4978_ (.A1(_0387_),
    .A2(_0401_),
    .ZN(_0402_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4979_ (.A1(_4273_),
    .A2(\as2650.cycle[1] ),
    .ZN(_0403_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4980_ (.I(_0403_),
    .Z(_0404_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4981_ (.I(_0404_),
    .Z(_0405_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4982_ (.I(_0405_),
    .Z(_0406_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _4983_ (.A1(_0318_),
    .A2(_0406_),
    .A3(_0330_),
    .A4(_0328_),
    .ZN(_0407_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4984_ (.A1(_0333_),
    .A2(_4417_),
    .B(_0407_),
    .ZN(_0408_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4985_ (.A1(_4350_),
    .A2(_0303_),
    .A3(_0408_),
    .ZN(_0409_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4986_ (.I(_4414_),
    .Z(_0410_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4987_ (.I(_0410_),
    .Z(_0411_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4988_ (.I(_0411_),
    .Z(_0412_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4989_ (.I(_0412_),
    .Z(_0413_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4990_ (.I(_4442_),
    .Z(_0414_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4991_ (.I(_0414_),
    .Z(_0415_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _4992_ (.A1(_0413_),
    .A2(_4366_),
    .A3(_0358_),
    .A4(_0415_),
    .ZN(_0416_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _4993_ (.A1(_0384_),
    .A2(_0402_),
    .A3(_0409_),
    .A4(_0416_),
    .ZN(_0008_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4994_ (.I(_4409_),
    .Z(_0417_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4995_ (.I(_0417_),
    .Z(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4996_ (.A1(_0323_),
    .A2(_0403_),
    .ZN(_0419_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4997_ (.A1(_0419_),
    .A2(_0325_),
    .ZN(_0420_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4998_ (.A1(_0413_),
    .A2(_0418_),
    .B1(_0420_),
    .B2(_4432_),
    .ZN(_0421_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4999_ (.A1(\as2650.cycle[2] ),
    .A2(_0296_),
    .ZN(_0422_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5000_ (.A1(_4351_),
    .A2(_0421_),
    .B(_0422_),
    .ZN(_0006_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5001_ (.I(_4367_),
    .Z(_0423_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5002_ (.I(_0423_),
    .Z(_0424_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5003_ (.I(_4324_),
    .Z(_0425_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5004_ (.I(_0365_),
    .Z(_0426_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _5005_ (.A1(_0424_),
    .A2(_0425_),
    .A3(_0298_),
    .A4(_0426_),
    .ZN(_0427_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5006_ (.A1(_0313_),
    .A2(_0294_),
    .B(_0427_),
    .ZN(_0005_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5007_ (.I(_4294_),
    .Z(_0428_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5008_ (.I(_4296_),
    .Z(_0429_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5009_ (.A1(_0428_),
    .A2(_0429_),
    .ZN(_0430_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5010_ (.A1(\as2650.cycle[3] ),
    .A2(_0296_),
    .ZN(_0431_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5011_ (.A1(_0366_),
    .A2(_0430_),
    .B(_0431_),
    .ZN(_0007_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5012_ (.I(_4290_),
    .Z(_0432_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5013_ (.I(_0432_),
    .Z(_0433_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5014_ (.I(_4288_),
    .Z(_0434_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5015_ (.I(_0434_),
    .Z(_0435_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5016_ (.I(_0435_),
    .Z(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5017_ (.I(_0429_),
    .Z(_0437_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5018_ (.I(_4242_),
    .Z(_0438_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _5019_ (.A1(_0437_),
    .A2(_0394_),
    .A3(_0438_),
    .A4(_0300_),
    .ZN(_0439_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5020_ (.A1(_0357_),
    .A2(_4442_),
    .ZN(_0440_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5021_ (.I(_0440_),
    .Z(_0441_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5022_ (.I(_4281_),
    .Z(_0442_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5023_ (.A1(_4280_),
    .A2(_4285_),
    .ZN(_0443_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _5024_ (.A1(_0438_),
    .A2(_0442_),
    .A3(_0443_),
    .B1(_4266_),
    .B2(_4275_),
    .ZN(_0444_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5025_ (.I(_4325_),
    .Z(_0445_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5026_ (.A1(_4313_),
    .A2(_0445_),
    .ZN(_0446_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _5027_ (.A1(_4277_),
    .A2(_4381_),
    .A3(_4056_),
    .ZN(_0447_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5028_ (.I(_0447_),
    .Z(_0448_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5029_ (.A1(_0448_),
    .A2(_4317_),
    .ZN(_0449_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5030_ (.A1(_4437_),
    .A2(_0381_),
    .B1(_0446_),
    .B2(_0449_),
    .ZN(_0450_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5031_ (.A1(_0383_),
    .A2(_4370_),
    .A3(_0303_),
    .ZN(_0451_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5032_ (.A1(_0353_),
    .A2(_4349_),
    .B(_0320_),
    .ZN(_0452_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5033_ (.A1(_0451_),
    .A2(_0452_),
    .ZN(_0453_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5034_ (.I(_4320_),
    .Z(_0454_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5035_ (.A1(_0299_),
    .A2(_0453_),
    .B1(_0446_),
    .B2(_0454_),
    .ZN(_0455_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5036_ (.A1(_4371_),
    .A2(_0450_),
    .B(_0455_),
    .ZN(_0456_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _5037_ (.A1(_0436_),
    .A2(_0439_),
    .B1(_0441_),
    .B2(_0444_),
    .C(_0456_),
    .ZN(_0457_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5038_ (.I(_0339_),
    .Z(_0458_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5039_ (.A1(_0413_),
    .A2(_0300_),
    .B(_0415_),
    .ZN(_0459_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _5040_ (.I(\as2650.addr_buff[7] ),
    .ZN(_0460_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5041_ (.I(_0460_),
    .Z(_0461_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5042_ (.A1(\as2650.cycle[13] ),
    .A2(_4447_),
    .ZN(_0462_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5043_ (.I(_0462_),
    .Z(_0463_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5044_ (.A1(_0461_),
    .A2(_0463_),
    .ZN(_0464_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5045_ (.I(_0432_),
    .Z(_0465_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5046_ (.I(_4242_),
    .Z(_0466_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5047_ (.A1(_0436_),
    .A2(_0464_),
    .B(_0465_),
    .C(_0466_),
    .ZN(_0467_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5048_ (.I(_4259_),
    .Z(_0468_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5049_ (.I(_0468_),
    .Z(_0469_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _5050_ (.A1(_0433_),
    .A2(_0458_),
    .B1(_0459_),
    .B2(_0467_),
    .C(_0469_),
    .ZN(_0470_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5051_ (.A1(_0428_),
    .A2(_4222_),
    .ZN(_0471_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5052_ (.I(_4085_),
    .Z(_0472_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5053_ (.I(_4396_),
    .Z(_0473_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5054_ (.A1(_4381_),
    .A2(_4234_),
    .ZN(_0474_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _5055_ (.A1(_0472_),
    .A2(_0473_),
    .A3(_0474_),
    .ZN(_0475_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5056_ (.I(_4086_),
    .Z(_0476_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5057_ (.A1(_4060_),
    .A2(_0476_),
    .ZN(_0477_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5058_ (.A1(_4386_),
    .A2(_0371_),
    .ZN(_0478_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _5059_ (.A1(_0477_),
    .A2(_4379_),
    .A3(_0478_),
    .ZN(_0479_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5060_ (.A1(_4372_),
    .A2(_0472_),
    .ZN(_0480_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5061_ (.I(_4378_),
    .Z(_0481_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5062_ (.A1(_4386_),
    .A2(_4382_),
    .ZN(_0482_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _5063_ (.A1(_0480_),
    .A2(_0481_),
    .A3(_0482_),
    .ZN(_0483_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5064_ (.A1(_0479_),
    .A2(_0483_),
    .ZN(_0484_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5065_ (.A1(_0475_),
    .A2(_0484_),
    .ZN(_0485_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _5066_ (.A1(_4387_),
    .A2(_4248_),
    .A3(_0473_),
    .A4(_4382_),
    .ZN(_0486_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5067_ (.A1(_4384_),
    .A2(_0486_),
    .ZN(_0487_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5068_ (.A1(_4398_),
    .A2(_0478_),
    .ZN(_0488_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5069_ (.I(_0488_),
    .Z(_0489_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5070_ (.I(_4391_),
    .Z(_0490_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5071_ (.I(_0481_),
    .Z(_0491_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5072_ (.I(_4079_),
    .Z(_0492_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5073_ (.I(_0492_),
    .Z(_0493_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5074_ (.I(_4055_),
    .Z(_0494_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5075_ (.A1(_0494_),
    .A2(_4419_),
    .ZN(_0495_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5076_ (.I(_0495_),
    .Z(_0496_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5077_ (.A1(_0493_),
    .A2(_0496_),
    .B(_4230_),
    .ZN(_0497_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _5078_ (.A1(_0305_),
    .A2(_0490_),
    .A3(_0491_),
    .A4(_0497_),
    .ZN(_0498_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _5079_ (.A1(_0485_),
    .A2(_0487_),
    .A3(_0489_),
    .A4(_0498_),
    .ZN(_0499_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5080_ (.A1(_0471_),
    .A2(_0499_),
    .B(_0433_),
    .ZN(_0500_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _5081_ (.A1(_4297_),
    .A2(_4094_),
    .A3(_0473_),
    .A4(_4382_),
    .ZN(_0501_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5082_ (.I(_0501_),
    .Z(_0502_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5083_ (.I(_0502_),
    .Z(_0503_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _5084_ (.A1(_4236_),
    .A2(_4257_),
    .B1(_4446_),
    .B2(_0503_),
    .C(_4312_),
    .ZN(_0504_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5085_ (.A1(_0500_),
    .A2(_0504_),
    .B(_4363_),
    .ZN(_0505_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5086_ (.A1(_0433_),
    .A2(_0457_),
    .B(_0470_),
    .C(_0505_),
    .ZN(_0000_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5087_ (.I(net27),
    .ZN(net14));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5088_ (.I(\as2650.r123[3][0] ),
    .Z(_0506_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5089_ (.I(_0506_),
    .Z(_0014_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5090_ (.I(\as2650.r123[3][1] ),
    .Z(_0507_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5091_ (.I(_0507_),
    .Z(_0015_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5092_ (.I(\as2650.r123[3][2] ),
    .Z(_0508_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5093_ (.I(_0508_),
    .Z(_0016_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5094_ (.I(\as2650.r123[3][3] ),
    .Z(_0509_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5095_ (.I(_0509_),
    .Z(_0017_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5096_ (.I(\as2650.r123[3][4] ),
    .Z(_0510_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5097_ (.I(_0510_),
    .Z(_0018_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5098_ (.I(\as2650.r123[3][5] ),
    .Z(_0511_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5099_ (.I(_0511_),
    .Z(_0019_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5100_ (.I(\as2650.r123[3][6] ),
    .Z(_0512_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5101_ (.I(_0512_),
    .Z(_0020_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5102_ (.I(\as2650.r123[3][7] ),
    .Z(_0513_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5103_ (.I(_0513_),
    .Z(_0021_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5104_ (.I(\as2650.r123[0][0] ),
    .ZN(_0514_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5105_ (.A1(\as2650.cycle[0] ),
    .A2(\as2650.cycle[8] ),
    .ZN(_0515_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5106_ (.A1(_4309_),
    .A2(_0515_),
    .ZN(_0516_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5107_ (.A1(_4064_),
    .A2(_0516_),
    .ZN(_0517_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5108_ (.A1(_4356_),
    .A2(_0517_),
    .ZN(_0518_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5109_ (.A1(_4393_),
    .A2(_0518_),
    .ZN(_0519_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5110_ (.A1(_0370_),
    .A2(_4305_),
    .ZN(_0520_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _5111_ (.A1(_4438_),
    .A2(_0519_),
    .A3(_0520_),
    .ZN(_0521_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5112_ (.I(_0521_),
    .Z(_0522_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5113_ (.I(_0522_),
    .Z(_0523_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5114_ (.I(_4064_),
    .Z(_0524_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _5115_ (.A1(_0524_),
    .A2(\as2650.cycle[0] ),
    .A3(_0492_),
    .A4(_4245_),
    .ZN(_0525_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5116_ (.I(_0525_),
    .Z(_0526_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5117_ (.A1(_4045_),
    .A2(_4261_),
    .ZN(_0527_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _5118_ (.A1(_4347_),
    .A2(_4333_),
    .A3(_0527_),
    .ZN(_0528_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5119_ (.A1(\as2650.cycle[5] ),
    .A2(\as2650.cycle[4] ),
    .ZN(_0529_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5120_ (.A1(_4386_),
    .A2(\as2650.cycle[8] ),
    .ZN(_0530_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5121_ (.A1(_0529_),
    .A2(_0530_),
    .ZN(_0531_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5122_ (.I(\as2650.addr_buff[6] ),
    .Z(_0532_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5123_ (.I(\as2650.addr_buff[5] ),
    .Z(_0533_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5124_ (.A1(_0532_),
    .A2(_0533_),
    .ZN(_0534_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5125_ (.A1(_0531_),
    .A2(_0534_),
    .ZN(_0535_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5126_ (.A1(_0528_),
    .A2(_0535_),
    .Z(_0536_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5127_ (.A1(_4413_),
    .A2(_0526_),
    .A3(_0536_),
    .ZN(_0537_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _5128_ (.A1(_0529_),
    .A2(_0323_),
    .A3(_0525_),
    .Z(_0538_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5129_ (.A1(\as2650.idx_ctrl[1] ),
    .A2(\as2650.idx_ctrl[0] ),
    .Z(_0539_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5130_ (.I(_0539_),
    .Z(_0540_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5131_ (.I(_0540_),
    .Z(_0541_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5132_ (.I(_0541_),
    .Z(_0542_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _5133_ (.A1(_4338_),
    .A2(_0542_),
    .A3(_0530_),
    .Z(_0543_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _5134_ (.A1(_0317_),
    .A2(_0528_),
    .A3(_0538_),
    .A4(_0543_),
    .ZN(_0544_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _5135_ (.A1(_0368_),
    .A2(_0302_),
    .A3(_0519_),
    .Z(_0545_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5136_ (.A1(_4438_),
    .A2(_0447_),
    .ZN(_0546_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5137_ (.I(_0518_),
    .Z(_0547_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _5138_ (.A1(_4449_),
    .A2(_0493_),
    .A3(_0546_),
    .A4(_0547_),
    .ZN(_0548_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5139_ (.I(_4082_),
    .Z(_0549_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5140_ (.I(_0515_),
    .Z(_0550_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _5141_ (.A1(_0549_),
    .A2(_4310_),
    .A3(_0550_),
    .ZN(_0551_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5142_ (.A1(\as2650.cycle[6] ),
    .A2(_4260_),
    .ZN(_0552_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _5143_ (.A1(_4373_),
    .A2(_4319_),
    .A3(_0552_),
    .ZN(_0553_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5144_ (.A1(_0551_),
    .A2(_0553_),
    .ZN(_0554_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5145_ (.I(_0524_),
    .Z(_0555_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5146_ (.I(_0550_),
    .Z(_0556_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5147_ (.A1(_4046_),
    .A2(_4438_),
    .ZN(_0557_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5148_ (.A1(_4057_),
    .A2(_0492_),
    .ZN(_0558_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _5149_ (.A1(_4310_),
    .A2(_0556_),
    .A3(_0557_),
    .A4(_0558_),
    .ZN(_0559_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5150_ (.I(_0517_),
    .Z(_0560_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5151_ (.A1(_4356_),
    .A2(_4344_),
    .ZN(_0561_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5152_ (.I(_0561_),
    .Z(_0562_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5153_ (.A1(_4282_),
    .A2(_0492_),
    .A3(_0542_),
    .ZN(_0563_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5154_ (.A1(_4297_),
    .A2(_0473_),
    .ZN(_0564_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _5155_ (.A1(_4170_),
    .A2(_0562_),
    .A3(_0563_),
    .A4(_0564_),
    .ZN(_0565_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5156_ (.I(_0565_),
    .ZN(_0566_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5157_ (.A1(_0560_),
    .A2(_0566_),
    .ZN(_0567_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5158_ (.A1(_0555_),
    .A2(_0559_),
    .B(_0567_),
    .ZN(_0568_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _5159_ (.A1(_0545_),
    .A2(_0548_),
    .A3(_0554_),
    .A4(_0568_),
    .ZN(_0569_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _5160_ (.A1(_0523_),
    .A2(_0537_),
    .A3(_0544_),
    .A4(_0569_),
    .Z(_0570_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5161_ (.A1(_0477_),
    .A2(_0570_),
    .ZN(_0571_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _5162_ (.A1(_0477_),
    .A2(_0491_),
    .A3(_0482_),
    .ZN(_0572_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5163_ (.A1(_0488_),
    .A2(_0572_),
    .ZN(_0573_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5164_ (.I(_0573_),
    .Z(_0574_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5165_ (.A1(_0547_),
    .A2(_0574_),
    .ZN(_0575_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _5166_ (.A1(_4259_),
    .A2(_0571_),
    .A3(_0575_),
    .ZN(_0576_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5167_ (.I(_0576_),
    .Z(_0577_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5168_ (.I(_0577_),
    .Z(_0578_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5169_ (.I(_0571_),
    .Z(_0579_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5170_ (.I(_0567_),
    .Z(_0580_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5171_ (.A1(_4389_),
    .A2(_4299_),
    .ZN(_0581_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _5172_ (.A1(_4230_),
    .A2(_0496_),
    .A3(_0581_),
    .ZN(_0582_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5173_ (.I(_0582_),
    .Z(_0583_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _5174_ (.I(\as2650.holding_reg[0] ),
    .ZN(_0584_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5175_ (.I(_4394_),
    .Z(_0585_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5176_ (.I0(_0584_),
    .I1(_4164_),
    .S(_0585_),
    .Z(_0586_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5177_ (.I(_0539_),
    .Z(_0587_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5178_ (.I(_4160_),
    .Z(_0588_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5179_ (.I(_0588_),
    .Z(_0589_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5180_ (.A1(_0589_),
    .A2(_0539_),
    .ZN(_0590_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5181_ (.I(_4375_),
    .Z(_0591_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _5182_ (.A1(_4164_),
    .A2(_0587_),
    .B(_0590_),
    .C(_0591_),
    .ZN(_0592_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5183_ (.A1(_0584_),
    .A2(_4395_),
    .ZN(_0593_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5184_ (.A1(_0586_),
    .A2(_0592_),
    .A3(_0593_),
    .ZN(_0594_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5185_ (.I(_0591_),
    .Z(_0595_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5186_ (.I(\as2650.idx_ctrl[1] ),
    .Z(_0596_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5187_ (.I(\as2650.idx_ctrl[0] ),
    .Z(_0597_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5188_ (.A1(_0596_),
    .A2(_0597_),
    .ZN(_0598_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5189_ (.I(_0598_),
    .Z(_0599_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5190_ (.A1(_4193_),
    .A2(_0599_),
    .Z(_0600_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5191_ (.I(_0589_),
    .Z(_0601_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5192_ (.I(_0591_),
    .Z(_0602_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5193_ (.A1(_0601_),
    .A2(_0599_),
    .B(_0602_),
    .ZN(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5194_ (.A1(\as2650.holding_reg[0] ),
    .A2(_0591_),
    .ZN(_0604_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5195_ (.A1(_4193_),
    .A2(_4376_),
    .B(_0604_),
    .ZN(_0605_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _5196_ (.A1(_0584_),
    .A2(_0595_),
    .B1(_0600_),
    .B2(_0603_),
    .C(_0605_),
    .ZN(_0606_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5197_ (.A1(_0594_),
    .A2(_0606_),
    .Z(_0607_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5198_ (.I(_0607_),
    .Z(_0608_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5199_ (.I(\as2650.psl[3] ),
    .Z(_0609_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5200_ (.I(\as2650.carry ),
    .Z(_0610_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5201_ (.A1(_0609_),
    .A2(_0610_),
    .ZN(_0611_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5202_ (.I(_0611_),
    .Z(_0612_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5203_ (.A1(_0608_),
    .A2(_0612_),
    .Z(_0613_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5204_ (.I(_4389_),
    .ZN(_0614_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5205_ (.I(_0614_),
    .Z(_0615_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5206_ (.A1(_0615_),
    .A2(_4251_),
    .ZN(_0616_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5207_ (.A1(_0608_),
    .A2(_0612_),
    .B(_0616_),
    .ZN(_0617_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5208_ (.I(\as2650.carry ),
    .ZN(_0618_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5209_ (.A1(\as2650.psl[3] ),
    .A2(_0618_),
    .ZN(_0619_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5210_ (.A1(_0614_),
    .A2(_4230_),
    .ZN(_0620_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5211_ (.I(_0620_),
    .Z(_0621_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5212_ (.A1(_0607_),
    .A2(_0619_),
    .B(_0621_),
    .ZN(_0622_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5213_ (.A1(_0608_),
    .A2(_0619_),
    .B(_0622_),
    .ZN(_0623_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5214_ (.A1(_4390_),
    .A2(_0495_),
    .ZN(_0624_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5215_ (.I(_0624_),
    .Z(_0625_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _5216_ (.I(_0625_),
    .ZN(_0626_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5217_ (.A1(_0605_),
    .A2(_0592_),
    .A3(_0593_),
    .ZN(_0627_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5218_ (.I(_0581_),
    .Z(_0628_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5219_ (.A1(_0592_),
    .A2(_0593_),
    .B(_0605_),
    .ZN(_0629_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5220_ (.I(_0370_),
    .Z(_0630_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5221_ (.A1(_4303_),
    .A2(_0630_),
    .ZN(_0631_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5222_ (.A1(_4390_),
    .A2(_0631_),
    .ZN(_0632_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5223_ (.A1(_0629_),
    .A2(_0632_),
    .Z(_0633_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _5224_ (.A1(_0626_),
    .A2(_0627_),
    .B1(_0607_),
    .B2(_0628_),
    .C(_0633_),
    .ZN(_0634_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _5225_ (.A1(_0613_),
    .A2(_0617_),
    .B(_0623_),
    .C(_0634_),
    .ZN(_0635_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5226_ (.I(_0582_),
    .Z(_0636_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5227_ (.A1(_0636_),
    .A2(_0605_),
    .ZN(_0637_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _5228_ (.A1(_0583_),
    .A2(_0635_),
    .B(_0637_),
    .ZN(_0638_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5229_ (.A1(_0330_),
    .A2(_0325_),
    .ZN(_0639_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5230_ (.I(_0599_),
    .Z(_0640_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5231_ (.I(_0640_),
    .Z(_0641_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _5232_ (.A1(_0314_),
    .A2(_0639_),
    .A3(_0641_),
    .A4(_0531_),
    .ZN(_0642_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _5233_ (.A1(_0318_),
    .A2(_0526_),
    .A3(_0528_),
    .A4(_0642_),
    .ZN(_0643_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5234_ (.I(_0643_),
    .Z(_0644_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5235_ (.I(_0596_),
    .ZN(_0645_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5236_ (.A1(_0645_),
    .A2(_0597_),
    .ZN(_0646_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5237_ (.I(\as2650.idx_ctrl[0] ),
    .ZN(_0647_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5238_ (.A1(_0596_),
    .A2(_0647_),
    .ZN(_0648_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5239_ (.A1(_0646_),
    .A2(_0648_),
    .ZN(_0649_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5240_ (.A1(_4193_),
    .A2(_0649_),
    .Z(_0650_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5241_ (.I(_0650_),
    .Z(_0651_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5242_ (.I(_0537_),
    .Z(_0652_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5243_ (.I(\as2650.addr_buff[5] ),
    .ZN(_0653_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5244_ (.A1(_0532_),
    .A2(_0653_),
    .ZN(_0654_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5245_ (.I(_0654_),
    .Z(_0655_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5246_ (.I(_0532_),
    .ZN(_0656_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5247_ (.A1(_0656_),
    .A2(_0533_),
    .ZN(_0657_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5248_ (.A1(_0655_),
    .A2(_0657_),
    .ZN(_0658_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5249_ (.A1(_4165_),
    .A2(_0658_),
    .Z(_0659_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5250_ (.I(_0659_),
    .Z(_0660_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5251_ (.I(_0537_),
    .Z(_0661_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5252_ (.I(_0601_),
    .Z(_0662_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5253_ (.I(_0662_),
    .Z(_0663_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5254_ (.I(_0545_),
    .Z(_0664_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5255_ (.A1(_0663_),
    .A2(_0664_),
    .ZN(_0665_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5256_ (.I(_0630_),
    .Z(_0666_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5257_ (.A1(_0666_),
    .A2(_4307_),
    .A3(_0519_),
    .ZN(_0667_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5258_ (.I(_0667_),
    .Z(_0668_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5259_ (.I(_0668_),
    .Z(_0669_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _5260_ (.A1(_4069_),
    .A2(_4074_),
    .A3(_4080_),
    .Z(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5261_ (.I(_0670_),
    .Z(_0671_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5262_ (.I(_0671_),
    .Z(_0672_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5263_ (.A1(_0609_),
    .A2(_0672_),
    .B(_0612_),
    .ZN(_0673_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5264_ (.I(_4209_),
    .Z(_0674_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5265_ (.I(net7),
    .Z(_0675_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5266_ (.I(_0675_),
    .Z(_0676_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5267_ (.A1(_0370_),
    .A2(_4326_),
    .ZN(_0677_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5268_ (.A1(_4322_),
    .A2(_0677_),
    .ZN(_0678_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5269_ (.A1(_4045_),
    .A2(_4344_),
    .ZN(_0679_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5270_ (.A1(_4393_),
    .A2(_0678_),
    .A3(_0679_),
    .ZN(_0680_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5271_ (.A1(_0560_),
    .A2(_0680_),
    .ZN(_0681_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5272_ (.I(_0681_),
    .Z(_0682_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5273_ (.I(_0681_),
    .Z(_0683_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5274_ (.A1(_4216_),
    .A2(_0683_),
    .ZN(_0684_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5275_ (.I(_0521_),
    .Z(_0685_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5276_ (.A1(_0676_),
    .A2(_0682_),
    .B(_0684_),
    .C(_0685_),
    .ZN(_0686_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5277_ (.A1(_0674_),
    .A2(_0522_),
    .B(_0686_),
    .C(_0668_),
    .ZN(_0687_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5278_ (.A1(_0367_),
    .A2(_0302_),
    .A3(_0519_),
    .ZN(_0688_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5279_ (.I(_0688_),
    .Z(_0689_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5280_ (.A1(_0669_),
    .A2(_0673_),
    .B(_0687_),
    .C(_0689_),
    .ZN(_0690_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5281_ (.A1(_0661_),
    .A2(_0665_),
    .A3(_0690_),
    .ZN(_0691_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5282_ (.I(_0544_),
    .Z(_0692_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5283_ (.A1(_0652_),
    .A2(_0660_),
    .B(_0691_),
    .C(_0692_),
    .ZN(_0693_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5284_ (.I(_0567_),
    .Z(_0694_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5285_ (.A1(_0644_),
    .A2(_0651_),
    .B(_0693_),
    .C(_0694_),
    .ZN(_0695_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5286_ (.A1(_0580_),
    .A2(_0638_),
    .B(_0695_),
    .ZN(_0696_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5287_ (.I(_0696_),
    .ZN(_0697_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5288_ (.I(_0663_),
    .Z(_0698_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5289_ (.I(\as2650.psu[0] ),
    .Z(_0699_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5290_ (.I(_0699_),
    .Z(_0700_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5291_ (.I(\as2650.psu[1] ),
    .ZN(_0701_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5292_ (.I(_0701_),
    .Z(_0702_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5293_ (.A1(_0700_),
    .A2(_0702_),
    .ZN(_0703_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5294_ (.I(_0703_),
    .Z(_0704_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5295_ (.I(_0704_),
    .Z(_0705_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5296_ (.I(\as2650.psu[0] ),
    .ZN(_0706_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5297_ (.I(_0706_),
    .Z(_0707_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5298_ (.I(\as2650.psu[1] ),
    .Z(_0708_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5299_ (.A1(_0707_),
    .A2(_0708_),
    .ZN(_0709_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5300_ (.I(_0709_),
    .Z(_0710_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5301_ (.I(_0710_),
    .Z(_0711_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5302_ (.A1(\as2650.psu[0] ),
    .A2(\as2650.psu[1] ),
    .ZN(_0712_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5303_ (.I(_0712_),
    .Z(_0713_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5304_ (.I(_0713_),
    .Z(_0714_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5305_ (.I(_0714_),
    .Z(_0715_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _5306_ (.A1(\as2650.stack[5][8] ),
    .A2(_0705_),
    .B1(_0711_),
    .B2(\as2650.stack[4][8] ),
    .C1(\as2650.stack[7][8] ),
    .C2(_0715_),
    .ZN(_0716_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5307_ (.A1(_0707_),
    .A2(_0702_),
    .ZN(_0717_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5308_ (.I(_0717_),
    .Z(_0718_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5309_ (.I(_0718_),
    .Z(_0719_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5310_ (.I(\as2650.psu[2] ),
    .ZN(_0720_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5311_ (.A1(_0720_),
    .A2(_0712_),
    .Z(_0721_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5312_ (.I(_0721_),
    .Z(_0722_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5313_ (.I(_0722_),
    .Z(_0723_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5314_ (.A1(\as2650.stack[6][8] ),
    .A2(_0719_),
    .B(_0723_),
    .ZN(_0724_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5315_ (.I(_0703_),
    .Z(_0725_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5316_ (.I(_0709_),
    .Z(_0726_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5317_ (.A1(\as2650.stack[1][8] ),
    .A2(_0725_),
    .B1(_0726_),
    .B2(\as2650.stack[0][8] ),
    .ZN(_0727_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5318_ (.I(_0727_),
    .ZN(_0728_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _5319_ (.A1(\as2650.stack[3][8] ),
    .A2(_0715_),
    .B1(_0719_),
    .B2(\as2650.stack[2][8] ),
    .C(_0728_),
    .ZN(_0729_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _5320_ (.A1(_0716_),
    .A2(_0724_),
    .B1(_0729_),
    .B2(_0723_),
    .ZN(_0730_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5321_ (.A1(_4380_),
    .A2(_0474_),
    .ZN(_0731_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5322_ (.I(_0731_),
    .Z(_0732_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5323_ (.I(_0732_),
    .Z(_0733_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5324_ (.A1(_0733_),
    .A2(_0547_),
    .ZN(_0734_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5325_ (.I0(_0698_),
    .I1(_0730_),
    .S(_0734_),
    .Z(_0735_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5326_ (.I(_4357_),
    .Z(_0736_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5327_ (.I(_0736_),
    .Z(_0737_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5328_ (.A1(_4398_),
    .A2(_0482_),
    .ZN(_0738_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5329_ (.I(_0738_),
    .Z(_0739_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5330_ (.A1(_0737_),
    .A2(_0739_),
    .ZN(_0740_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5331_ (.A1(_0551_),
    .A2(_0740_),
    .ZN(_0741_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5332_ (.A1(_0575_),
    .A2(_0741_),
    .ZN(_0742_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5333_ (.I(_0742_),
    .Z(_0743_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5334_ (.I(_0743_),
    .ZN(_0744_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5335_ (.I(_0576_),
    .Z(_0745_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _5336_ (.A1(_0579_),
    .A2(_0697_),
    .B1(_0735_),
    .B2(_0744_),
    .C(_0745_),
    .ZN(_0746_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5337_ (.A1(_0514_),
    .A2(_0578_),
    .B(_0746_),
    .ZN(_0022_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5338_ (.I(\as2650.r123[0][1] ),
    .ZN(_0747_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5339_ (.I(_0694_),
    .Z(_0748_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5340_ (.A1(\as2650.holding_reg[1] ),
    .A2(_4376_),
    .ZN(_0749_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5341_ (.A1(_4208_),
    .A2(_0602_),
    .B(_0749_),
    .ZN(_0750_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5342_ (.A1(_4147_),
    .A2(_4153_),
    .A3(_0598_),
    .ZN(_0751_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5343_ (.I(_4150_),
    .Z(_0752_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _5344_ (.I(_0752_),
    .ZN(_0753_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5345_ (.A1(_0753_),
    .A2(_0539_),
    .B(_4394_),
    .ZN(_0754_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5346_ (.A1(\as2650.holding_reg[1] ),
    .A2(_0585_),
    .B1(_0751_),
    .B2(_0754_),
    .ZN(_0755_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5347_ (.I(_0755_),
    .Z(_0756_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5348_ (.A1(_0750_),
    .A2(_0756_),
    .Z(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5349_ (.I(_0757_),
    .Z(_0758_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5350_ (.A1(_0607_),
    .A2(_0619_),
    .ZN(_0759_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5351_ (.A1(_0594_),
    .A2(_0759_),
    .ZN(_0760_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5352_ (.A1(_0758_),
    .A2(_0760_),
    .B(_0621_),
    .ZN(_0761_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5353_ (.A1(_0758_),
    .A2(_0760_),
    .B(_0761_),
    .ZN(_0762_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5354_ (.A1(_4148_),
    .A2(_4154_),
    .A3(_4394_),
    .ZN(_0763_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5355_ (.A1(\as2650.holding_reg[1] ),
    .A2(_0585_),
    .B(_0763_),
    .ZN(_0764_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5356_ (.A1(_0764_),
    .A2(_0755_),
    .Z(_0765_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5357_ (.A1(_0629_),
    .A2(_0611_),
    .B(_0627_),
    .ZN(_0766_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5358_ (.A1(_0765_),
    .A2(_0766_),
    .Z(_0767_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5359_ (.A1(_0765_),
    .A2(_0766_),
    .B(_4383_),
    .ZN(_0768_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5360_ (.A1(_0767_),
    .A2(_0768_),
    .ZN(_0769_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5361_ (.I(_0628_),
    .Z(_0770_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5362_ (.A1(_0764_),
    .A2(_0756_),
    .ZN(_0771_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5363_ (.A1(_0764_),
    .A2(_0756_),
    .ZN(_0772_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5364_ (.A1(_4391_),
    .A2(_0771_),
    .B(_0772_),
    .C(_0631_),
    .ZN(_0773_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5365_ (.A1(_0770_),
    .A2(_0758_),
    .B(_0773_),
    .C(_0636_),
    .ZN(_0774_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _5366_ (.A1(_0762_),
    .A2(_0769_),
    .A3(_0774_),
    .B1(_0750_),
    .B2(_0583_),
    .ZN(_0775_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5367_ (.I(_0752_),
    .Z(_0776_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5368_ (.I(_0776_),
    .Z(_0777_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5369_ (.I(_0777_),
    .Z(_0778_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5370_ (.I(_0545_),
    .Z(_0779_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _5371_ (.A1(_4413_),
    .A2(_0526_),
    .A3(_0536_),
    .Z(_0780_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5372_ (.I(_0780_),
    .Z(_0781_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5373_ (.I(_4215_),
    .Z(_0782_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5374_ (.I(_0548_),
    .Z(_0783_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5375_ (.I(net8),
    .Z(_0784_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5376_ (.I(_0784_),
    .Z(_0785_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5377_ (.I(_0785_),
    .Z(_0786_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5378_ (.I(_0786_),
    .Z(_0787_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5379_ (.I(_0682_),
    .Z(_0788_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5380_ (.A1(_4218_),
    .A2(_0788_),
    .ZN(_0789_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5381_ (.A1(_0787_),
    .A2(_0788_),
    .B(_0789_),
    .C(_0523_),
    .ZN(_0790_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5382_ (.I(_4144_),
    .Z(_0791_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5383_ (.A1(_4419_),
    .A2(_0447_),
    .ZN(_0792_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5384_ (.I(_0792_),
    .Z(_0793_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _5385_ (.A1(_0428_),
    .A2(_0493_),
    .A3(_0547_),
    .A4(_0793_),
    .ZN(_0794_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5386_ (.A1(_0791_),
    .A2(_0794_),
    .B(_0783_),
    .ZN(_0795_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _5387_ (.A1(_0782_),
    .A2(_0783_),
    .B1(_0790_),
    .B2(_0795_),
    .C(_0664_),
    .ZN(_0796_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5388_ (.A1(_0778_),
    .A2(_0779_),
    .B(_0781_),
    .C(_0796_),
    .ZN(_0797_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5389_ (.I(_4163_),
    .Z(_0798_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5390_ (.A1(\as2650.addr_buff[6] ),
    .A2(_0653_),
    .ZN(_0799_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5391_ (.A1(_0798_),
    .A2(_0654_),
    .B(_0799_),
    .ZN(_0800_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _5392_ (.A1(_4208_),
    .A2(_0798_),
    .A3(_0800_),
    .Z(_0801_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5393_ (.I(_0801_),
    .Z(_0802_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5394_ (.A1(_0652_),
    .A2(_0802_),
    .B(_0692_),
    .ZN(_0803_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5395_ (.A1(\as2650.idx_ctrl[1] ),
    .A2(_0647_),
    .ZN(_0804_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5396_ (.A1(_4176_),
    .A2(_0804_),
    .B(_0648_),
    .ZN(_0805_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _5397_ (.A1(_4208_),
    .A2(_0798_),
    .A3(_0805_),
    .Z(_0806_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5398_ (.I(_0806_),
    .ZN(_0807_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5399_ (.I(_0544_),
    .Z(_0808_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5400_ (.A1(_0797_),
    .A2(_0803_),
    .B1(_0807_),
    .B2(_0808_),
    .ZN(_0809_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5401_ (.A1(_0580_),
    .A2(_0809_),
    .ZN(_0810_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5402_ (.A1(_0748_),
    .A2(_0775_),
    .B(_0810_),
    .ZN(_0811_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5403_ (.I(_4358_),
    .Z(_0812_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5404_ (.I(_0812_),
    .Z(_0813_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5405_ (.I(_0813_),
    .Z(_0814_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5406_ (.I(_0488_),
    .Z(_0815_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5407_ (.A1(_0814_),
    .A2(_0815_),
    .A3(_0560_),
    .ZN(_0816_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5408_ (.I(_0816_),
    .Z(_0817_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5409_ (.I(_0817_),
    .Z(_0818_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5410_ (.A1(_0753_),
    .A2(_0818_),
    .ZN(_0819_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5411_ (.I(_0816_),
    .Z(_0820_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5412_ (.I(_0713_),
    .Z(_0821_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5413_ (.I(_0717_),
    .Z(_0822_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5414_ (.A1(\as2650.stack[7][9] ),
    .A2(_0821_),
    .B1(_0822_),
    .B2(\as2650.stack[6][9] ),
    .ZN(_0823_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5415_ (.I(_0703_),
    .Z(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5416_ (.I(_0721_),
    .Z(_0825_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _5417_ (.A1(\as2650.stack[5][9] ),
    .A2(_0824_),
    .B1(_0726_),
    .B2(\as2650.stack[4][9] ),
    .C(_0825_),
    .ZN(_0826_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5418_ (.I(_0709_),
    .Z(_0827_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5419_ (.A1(\as2650.stack[3][9] ),
    .A2(_0714_),
    .B1(_0704_),
    .B2(\as2650.stack[1][9] ),
    .ZN(_0828_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5420_ (.I(_0828_),
    .ZN(_0829_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _5421_ (.A1(\as2650.stack[0][9] ),
    .A2(_0827_),
    .B1(_0718_),
    .B2(\as2650.stack[2][9] ),
    .C(_0829_),
    .ZN(_0830_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5422_ (.I(_0722_),
    .Z(_0831_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _5423_ (.A1(_0823_),
    .A2(_0826_),
    .B1(_0830_),
    .B2(_0831_),
    .ZN(_0832_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5424_ (.A1(_0820_),
    .A2(_0832_),
    .ZN(_0833_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5425_ (.A1(_0743_),
    .A2(_0833_),
    .ZN(_0834_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _5426_ (.A1(_0571_),
    .A2(_0811_),
    .B1(_0819_),
    .B2(_0834_),
    .C(_0576_),
    .ZN(_0835_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5427_ (.A1(_0747_),
    .A2(_0578_),
    .B(_0835_),
    .ZN(_0023_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5428_ (.I(\as2650.r123[0][2] ),
    .ZN(_0836_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5429_ (.A1(\as2650.holding_reg[2] ),
    .A2(_0602_),
    .ZN(_0837_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5430_ (.A1(_4191_),
    .A2(_4377_),
    .B(_0837_),
    .ZN(_0838_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5431_ (.A1(_0636_),
    .A2(_0838_),
    .ZN(_0839_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5432_ (.I(_0585_),
    .Z(_0840_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5433_ (.A1(_4137_),
    .A2(_4142_),
    .A3(_4395_),
    .ZN(_0841_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5434_ (.A1(\as2650.holding_reg[2] ),
    .A2(_0840_),
    .B(_0841_),
    .ZN(_0842_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5435_ (.A1(_4137_),
    .A2(_4142_),
    .A3(_0599_),
    .ZN(_0843_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5436_ (.I(_4139_),
    .Z(_0844_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _5437_ (.I(_0844_),
    .ZN(_0845_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5438_ (.A1(_0845_),
    .A2(_0587_),
    .B(_4395_),
    .ZN(_0846_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _5439_ (.A1(\as2650.holding_reg[2] ),
    .A2(_0840_),
    .B1(_0843_),
    .B2(_0846_),
    .ZN(_0847_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5440_ (.A1(_0842_),
    .A2(_0847_),
    .ZN(_0848_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5441_ (.A1(_0842_),
    .A2(_0847_),
    .Z(_0849_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5442_ (.A1(_0848_),
    .A2(_0849_),
    .Z(_0850_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5443_ (.A1(_0771_),
    .A2(_0767_),
    .ZN(_0851_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5444_ (.A1(_0850_),
    .A2(_0851_),
    .Z(_0852_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5445_ (.I(_0849_),
    .Z(_0853_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5446_ (.I(_0850_),
    .Z(_0854_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5447_ (.A1(_4389_),
    .A2(_4299_),
    .Z(_0855_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _5448_ (.A1(_4251_),
    .A2(_0631_),
    .A3(_0855_),
    .ZN(_0856_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5449_ (.A1(_0624_),
    .A2(_0848_),
    .B(_0856_),
    .ZN(_0857_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _5450_ (.A1(_0632_),
    .A2(_0853_),
    .B1(_0854_),
    .B2(_0628_),
    .C(_0857_),
    .ZN(_0858_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _5451_ (.A1(_0586_),
    .A2(_0592_),
    .A3(_0593_),
    .Z(_0859_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5452_ (.A1(_0606_),
    .A2(_0619_),
    .B(_0859_),
    .ZN(_0860_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5453_ (.A1(_0750_),
    .A2(_0756_),
    .Z(_0861_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5454_ (.A1(_0765_),
    .A2(_0860_),
    .B(_0861_),
    .ZN(_0862_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5455_ (.A1(_0854_),
    .A2(_0862_),
    .B(_0621_),
    .ZN(_0863_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5456_ (.A1(_0854_),
    .A2(_0862_),
    .B(_0863_),
    .ZN(_0864_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5457_ (.A1(_4383_),
    .A2(_0852_),
    .B(_0858_),
    .C(_0864_),
    .ZN(_0865_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5458_ (.A1(_0839_),
    .A2(_0865_),
    .ZN(_0866_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5459_ (.A1(_4148_),
    .A2(_4154_),
    .B(_4164_),
    .ZN(_0867_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5460_ (.A1(_4191_),
    .A2(_0867_),
    .Z(_0868_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _5461_ (.A1(_4148_),
    .A2(_4154_),
    .A3(_4176_),
    .Z(_0869_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5462_ (.A1(_4190_),
    .A2(_0869_),
    .Z(_0870_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5463_ (.I(_0657_),
    .Z(_0871_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5464_ (.A1(_0654_),
    .A2(_0657_),
    .Z(_0872_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5465_ (.A1(_4143_),
    .A2(_0872_),
    .ZN(_0873_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _5466_ (.A1(_0655_),
    .A2(_0868_),
    .B1(_0870_),
    .B2(_0871_),
    .C(_0873_),
    .ZN(_0874_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5467_ (.I(_0874_),
    .ZN(_0875_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5468_ (.I(_0844_),
    .Z(_0876_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5469_ (.I(_0876_),
    .Z(_0877_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5470_ (.I(_0688_),
    .Z(_0878_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5471_ (.I(_0667_),
    .Z(_0879_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5472_ (.I(_4207_),
    .Z(_0880_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5473_ (.I(net9),
    .Z(_0881_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5474_ (.I(_0881_),
    .Z(_0882_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5475_ (.I(_0882_),
    .Z(_0883_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5476_ (.A1(_4214_),
    .A2(_0683_),
    .ZN(_0884_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5477_ (.A1(_0883_),
    .A2(_0682_),
    .B(_0884_),
    .C(_0685_),
    .ZN(_0885_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5478_ (.A1(_0880_),
    .A2(_0522_),
    .B(_0885_),
    .C(_0668_),
    .ZN(_0886_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5479_ (.A1(_4156_),
    .A2(_0879_),
    .B(_0886_),
    .ZN(_0887_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5480_ (.A1(_0878_),
    .A2(_0887_),
    .ZN(_0888_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5481_ (.A1(_0877_),
    .A2(_0878_),
    .B(_0661_),
    .C(_0888_),
    .ZN(_0889_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5482_ (.A1(_0652_),
    .A2(_0875_),
    .B(_0889_),
    .ZN(_0890_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5483_ (.A1(_0645_),
    .A2(_0597_),
    .ZN(_0891_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5484_ (.I(_0891_),
    .Z(_0892_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5485_ (.A1(_0892_),
    .A2(_0870_),
    .Z(_0893_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5486_ (.A1(_4143_),
    .A2(_0867_),
    .Z(_0894_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_4 _5487_ (.A1(_4144_),
    .A2(_0649_),
    .B1(_0894_),
    .B2(_0646_),
    .ZN(_0895_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5488_ (.A1(_0893_),
    .A2(_0895_),
    .ZN(_0896_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5489_ (.A1(_0528_),
    .A2(_0543_),
    .ZN(_0897_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _5490_ (.A1(_0318_),
    .A2(_0529_),
    .A3(_0324_),
    .A4(_0526_),
    .ZN(_0898_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5491_ (.A1(_0897_),
    .A2(_0898_),
    .ZN(_0899_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5492_ (.I0(_0890_),
    .I1(_0896_),
    .S(_0899_),
    .Z(_0900_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5493_ (.I0(_0866_),
    .I1(_0900_),
    .S(_0580_),
    .Z(_0901_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5494_ (.A1(\as2650.stack[7][10] ),
    .A2(_0821_),
    .B1(_0822_),
    .B2(\as2650.stack[6][10] ),
    .ZN(_0902_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _5495_ (.A1(\as2650.stack[5][10] ),
    .A2(_0725_),
    .B1(_0726_),
    .B2(\as2650.stack[4][10] ),
    .C(_0825_),
    .ZN(_0903_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5496_ (.A1(\as2650.stack[3][10] ),
    .A2(_0821_),
    .B1(_0822_),
    .B2(\as2650.stack[2][10] ),
    .ZN(_0904_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5497_ (.A1(\as2650.psu[2] ),
    .A2(_0713_),
    .Z(_0905_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5498_ (.I(_0905_),
    .Z(_0906_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _5499_ (.A1(\as2650.stack[1][10] ),
    .A2(_0824_),
    .B1(_0827_),
    .B2(\as2650.stack[0][10] ),
    .C(_0906_),
    .ZN(_0907_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _5500_ (.A1(_0902_),
    .A2(_0903_),
    .B1(_0904_),
    .B2(_0907_),
    .ZN(_0908_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5501_ (.A1(_0817_),
    .A2(_0908_),
    .ZN(_0909_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5502_ (.A1(_0845_),
    .A2(_0820_),
    .B(_0742_),
    .C(_0909_),
    .ZN(_0910_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5503_ (.A1(_0579_),
    .A2(_0901_),
    .B(_0910_),
    .C(_0577_),
    .ZN(_0911_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5504_ (.A1(_0836_),
    .A2(_0578_),
    .B(_0911_),
    .ZN(_0024_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5505_ (.I(\as2650.r123[0][3] ),
    .ZN(_0912_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5506_ (.I(_0567_),
    .Z(_0913_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5507_ (.I(_0856_),
    .Z(_0914_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5508_ (.A1(_4206_),
    .A2(_0595_),
    .ZN(_0915_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _5509_ (.A1(\as2650.holding_reg[3] ),
    .A2(_4377_),
    .B(_0915_),
    .ZN(_0916_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5510_ (.I(_0602_),
    .Z(_0917_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5511_ (.I(_4128_),
    .Z(_0918_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5512_ (.A1(_0918_),
    .A2(_0587_),
    .ZN(_0919_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5513_ (.A1(_4206_),
    .A2(_0540_),
    .B(_0919_),
    .C(_0595_),
    .ZN(_0920_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5514_ (.A1(\as2650.holding_reg[3] ),
    .A2(_0917_),
    .B(_0920_),
    .ZN(_0921_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5515_ (.A1(_0916_),
    .A2(_0921_),
    .Z(_0922_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5516_ (.A1(_0916_),
    .A2(_0921_),
    .ZN(_0923_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5517_ (.A1(_0922_),
    .A2(_0923_),
    .Z(_0924_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5518_ (.I(_0924_),
    .Z(_0925_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _5519_ (.A1(_0771_),
    .A2(_0767_),
    .A3(_0848_),
    .ZN(_0926_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5520_ (.A1(_0853_),
    .A2(_0926_),
    .B(_4383_),
    .ZN(_0927_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5521_ (.A1(_0770_),
    .A2(_0927_),
    .ZN(_0928_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5522_ (.A1(_0925_),
    .A2(_0928_),
    .ZN(_0929_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5523_ (.I(_0620_),
    .Z(_0930_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5524_ (.I(_0930_),
    .Z(_0931_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5525_ (.A1(_0838_),
    .A2(_0847_),
    .Z(_0932_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5526_ (.I(_0932_),
    .ZN(_0933_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _5527_ (.A1(_0850_),
    .A2(_0862_),
    .B(_0933_),
    .ZN(_0934_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5528_ (.A1(_0925_),
    .A2(_0934_),
    .Z(_0935_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _5529_ (.A1(_0616_),
    .A2(_0853_),
    .A3(_0925_),
    .A4(_0926_),
    .ZN(_0936_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5530_ (.A1(_0916_),
    .A2(_0921_),
    .Z(_0937_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _5531_ (.A1(_0626_),
    .A2(_0922_),
    .B1(_0937_),
    .B2(_0632_),
    .C(_0582_),
    .ZN(_0938_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _5532_ (.A1(_0931_),
    .A2(_0935_),
    .B(_0936_),
    .C(_0938_),
    .ZN(_0939_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _5533_ (.A1(_0914_),
    .A2(_0916_),
    .B1(_0929_),
    .B2(_0939_),
    .ZN(_0940_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5534_ (.I(_0804_),
    .Z(_0941_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _5535_ (.A1(_4136_),
    .A2(_4141_),
    .B1(_4147_),
    .B2(_4153_),
    .C(_0798_),
    .ZN(_0942_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5536_ (.A1(_4205_),
    .A2(_0942_),
    .Z(_0943_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5537_ (.A1(_0941_),
    .A2(_0943_),
    .Z(_0944_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5538_ (.A1(_4177_),
    .A2(_4178_),
    .ZN(_0945_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5539_ (.A1(_4191_),
    .A2(_0869_),
    .B(_4206_),
    .ZN(_0946_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _5540_ (.A1(_0945_),
    .A2(_0648_),
    .A3(_0946_),
    .B1(_0649_),
    .B2(_4134_),
    .ZN(_0947_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5541_ (.A1(_0944_),
    .A2(_0947_),
    .Z(_0948_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5542_ (.I(_0918_),
    .Z(_0949_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5543_ (.I(_4192_),
    .Z(_0950_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5544_ (.I(_4175_),
    .Z(_0951_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5545_ (.I(net10),
    .Z(_0952_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5546_ (.I(_0952_),
    .Z(_0953_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5547_ (.A1(_0953_),
    .A2(_0554_),
    .ZN(_0954_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5548_ (.A1(_4212_),
    .A2(_0554_),
    .B(_0954_),
    .C(_0521_),
    .ZN(_0955_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5549_ (.A1(_0951_),
    .A2(_0522_),
    .B(_0955_),
    .C(_0668_),
    .ZN(_0956_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5550_ (.A1(_0950_),
    .A2(_0879_),
    .B(_0956_),
    .C(_0689_),
    .ZN(_0957_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5551_ (.A1(_0949_),
    .A2(_0878_),
    .B(_0661_),
    .C(_0957_),
    .ZN(_0958_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5552_ (.I(_0658_),
    .Z(_0959_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5553_ (.A1(_0945_),
    .A2(_0799_),
    .A3(_0946_),
    .ZN(_0960_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _5554_ (.A1(_4207_),
    .A2(_0959_),
    .B1(_0943_),
    .B2(_0655_),
    .C(_0960_),
    .ZN(_0961_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5555_ (.I(_0961_),
    .Z(_0962_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5556_ (.A1(_0780_),
    .A2(_0962_),
    .ZN(_0963_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5557_ (.A1(_0958_),
    .A2(_0963_),
    .ZN(_0964_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5558_ (.A1(_0692_),
    .A2(_0964_),
    .ZN(_0965_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5559_ (.A1(_0808_),
    .A2(_0948_),
    .B(_0965_),
    .C(_0694_),
    .ZN(_0966_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5560_ (.A1(_0913_),
    .A2(_0940_),
    .B(_0966_),
    .ZN(_0967_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5561_ (.I(_0967_),
    .ZN(_0968_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5562_ (.I(_0949_),
    .Z(_0969_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _5563_ (.I(_0969_),
    .ZN(_0970_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5564_ (.A1(_0970_),
    .A2(_0818_),
    .ZN(_0971_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _5565_ (.A1(\as2650.stack[1][11] ),
    .A2(_0725_),
    .B1(_0726_),
    .B2(\as2650.stack[0][11] ),
    .C1(_0718_),
    .C2(\as2650.stack[2][11] ),
    .ZN(_0972_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5566_ (.I(_0905_),
    .Z(_0973_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5567_ (.A1(\as2650.stack[3][11] ),
    .A2(_0715_),
    .B(_0973_),
    .ZN(_0974_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _5568_ (.A1(\as2650.stack[5][11] ),
    .A2(_0704_),
    .B1(_0710_),
    .B2(\as2650.stack[4][11] ),
    .C1(\as2650.stack[7][11] ),
    .C2(_0713_),
    .ZN(_0975_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5569_ (.A1(_0906_),
    .A2(_0975_),
    .ZN(_0976_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5570_ (.A1(\as2650.stack[6][11] ),
    .A2(_0719_),
    .B(_0976_),
    .ZN(_0977_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _5571_ (.A1(_0972_),
    .A2(_0974_),
    .B(_0977_),
    .ZN(_0978_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5572_ (.A1(_0820_),
    .A2(_0978_),
    .ZN(_0979_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5573_ (.A1(_0743_),
    .A2(_0979_),
    .ZN(_0980_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _5574_ (.A1(_0571_),
    .A2(_0968_),
    .B1(_0971_),
    .B2(_0980_),
    .C(_0576_),
    .ZN(_0981_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5575_ (.A1(_0912_),
    .A2(_0578_),
    .B(_0981_),
    .ZN(_0025_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5576_ (.I(\as2650.r123[0][4] ),
    .ZN(_0982_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5577_ (.I(_0577_),
    .Z(_0983_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5578_ (.A1(_4175_),
    .A2(_4396_),
    .ZN(_0984_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5579_ (.A1(\as2650.holding_reg[4] ),
    .A2(_0917_),
    .ZN(_0985_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5580_ (.A1(_0984_),
    .A2(_0985_),
    .ZN(_0986_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5581_ (.A1(_0984_),
    .A2(_0985_),
    .Z(_0987_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5582_ (.I(_4118_),
    .Z(_0988_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5583_ (.A1(_0988_),
    .A2(_0540_),
    .ZN(_0989_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5584_ (.A1(_4125_),
    .A2(_0541_),
    .B(_0989_),
    .C(_4377_),
    .ZN(_0990_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5585_ (.A1(\as2650.holding_reg[4] ),
    .A2(_0917_),
    .B(_0990_),
    .ZN(_0991_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5586_ (.A1(_0987_),
    .A2(_0991_),
    .ZN(_0992_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5587_ (.I(_0992_),
    .ZN(_0993_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5588_ (.A1(_0987_),
    .A2(_0991_),
    .ZN(_0994_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5589_ (.A1(_0993_),
    .A2(_0994_),
    .ZN(_0995_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5590_ (.I(_0995_),
    .Z(_0996_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _5591_ (.A1(\as2650.holding_reg[3] ),
    .A2(_4378_),
    .B(_0915_),
    .C(_0921_),
    .ZN(_0997_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5592_ (.I(_0997_),
    .ZN(_0998_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5593_ (.A1(_0924_),
    .A2(_0934_),
    .B(_0998_),
    .ZN(_0999_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5594_ (.A1(_0996_),
    .A2(_0999_),
    .B(_0930_),
    .ZN(_1000_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5595_ (.A1(_0996_),
    .A2(_0999_),
    .B(_1000_),
    .ZN(_1001_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _5596_ (.A1(_0849_),
    .A2(_0937_),
    .A3(_0926_),
    .B(_0922_),
    .ZN(_1002_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5597_ (.A1(_0995_),
    .A2(_1002_),
    .Z(_1003_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5598_ (.I(_0616_),
    .Z(_1004_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5599_ (.A1(_0615_),
    .A2(_0496_),
    .ZN(_1005_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _5600_ (.A1(_0625_),
    .A2(_0992_),
    .B1(_0994_),
    .B2(_1005_),
    .C(_0856_),
    .ZN(_1006_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _5601_ (.A1(_0770_),
    .A2(_0996_),
    .B1(_1003_),
    .B2(_1004_),
    .C(_1006_),
    .ZN(_1007_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5602_ (.A1(_0636_),
    .A2(_0986_),
    .B1(_1001_),
    .B2(_1007_),
    .ZN(_1008_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5603_ (.I(_1008_),
    .Z(_1009_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5604_ (.A1(_0804_),
    .A2(_0891_),
    .ZN(_1010_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5605_ (.A1(_4133_),
    .A2(_0942_),
    .ZN(_1011_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5606_ (.A1(_4174_),
    .A2(_1011_),
    .Z(_1012_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5607_ (.A1(_4124_),
    .A2(_0945_),
    .Z(_1013_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _5608_ (.A1(_4125_),
    .A2(_1010_),
    .B1(_1012_),
    .B2(_0804_),
    .C1(_1013_),
    .C2(_0892_),
    .ZN(_1014_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5609_ (.I(_1014_),
    .Z(_1015_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5610_ (.I(_0780_),
    .Z(_1016_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5611_ (.I(_0988_),
    .Z(_1017_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5612_ (.I(_1017_),
    .Z(_1018_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5613_ (.I(net11),
    .Z(_1019_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5614_ (.I(_1019_),
    .Z(_1020_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5615_ (.I(_1020_),
    .Z(_1021_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5616_ (.I(_1021_),
    .Z(_1022_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5617_ (.I(_1022_),
    .Z(_1023_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5618_ (.I(_0683_),
    .Z(_1024_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5619_ (.A1(_4198_),
    .A2(_1024_),
    .ZN(_1025_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5620_ (.I(_0521_),
    .Z(_1026_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5621_ (.A1(_1023_),
    .A2(_0788_),
    .B(_1025_),
    .C(_1026_),
    .ZN(_1027_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5622_ (.I(_4202_),
    .Z(_1028_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5623_ (.A1(_1028_),
    .A2(_0794_),
    .B(_0548_),
    .ZN(_1029_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _5624_ (.A1(_0880_),
    .A2(_0783_),
    .B1(_1027_),
    .B2(_1029_),
    .C(_0664_),
    .ZN(_1030_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5625_ (.A1(_1018_),
    .A2(_0779_),
    .B(_1030_),
    .ZN(_1031_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5626_ (.I(_0655_),
    .Z(_1032_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5627_ (.A1(_0951_),
    .A2(_0872_),
    .ZN(_1033_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _5628_ (.A1(_1032_),
    .A2(_1012_),
    .B1(_1013_),
    .B2(_0871_),
    .C(_1033_),
    .ZN(_1034_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5629_ (.I(_1034_),
    .Z(_1035_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5630_ (.A1(_1016_),
    .A2(_1035_),
    .ZN(_1036_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5631_ (.A1(_1016_),
    .A2(_1031_),
    .B(_1036_),
    .C(_0808_),
    .ZN(_1037_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5632_ (.A1(_0644_),
    .A2(_1015_),
    .B(_1037_),
    .C(_0913_),
    .ZN(_1038_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5633_ (.A1(_0748_),
    .A2(_1009_),
    .B(_1038_),
    .ZN(_1039_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5634_ (.A1(\as2650.stack[3][12] ),
    .A2(_0714_),
    .B1(_0710_),
    .B2(\as2650.stack[0][12] ),
    .ZN(_1040_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5635_ (.I(_1040_),
    .ZN(_1041_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _5636_ (.A1(\as2650.stack[1][12] ),
    .A2(_0725_),
    .B1(_0822_),
    .B2(\as2650.stack[2][12] ),
    .C(_1041_),
    .ZN(_1042_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5637_ (.I(_0714_),
    .Z(_1043_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5638_ (.I(_0717_),
    .Z(_1044_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5639_ (.A1(\as2650.stack[7][12] ),
    .A2(_1043_),
    .B1(_1044_),
    .B2(\as2650.stack[6][12] ),
    .ZN(_1045_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5640_ (.I(_0721_),
    .Z(_1046_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5641_ (.I(_1046_),
    .Z(_1047_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _5642_ (.A1(\as2650.stack[5][12] ),
    .A2(_0824_),
    .B1(_0827_),
    .B2(\as2650.stack[4][12] ),
    .C(_1047_),
    .ZN(_1048_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _5643_ (.A1(_0831_),
    .A2(_1042_),
    .B1(_1045_),
    .B2(_1048_),
    .ZN(_1049_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5644_ (.A1(_0817_),
    .A2(_1049_),
    .ZN(_1050_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5645_ (.A1(_1018_),
    .A2(_0734_),
    .ZN(_1051_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5646_ (.A1(_0742_),
    .A2(_1050_),
    .A3(_1051_),
    .ZN(_1052_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5647_ (.A1(_0579_),
    .A2(_1039_),
    .B(_1052_),
    .C(_0745_),
    .ZN(_1053_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5648_ (.A1(_0982_),
    .A2(_0983_),
    .B(_1053_),
    .ZN(_0026_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5649_ (.I(\as2650.r123[0][5] ),
    .ZN(_1054_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5650_ (.I(_4116_),
    .Z(_1055_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5651_ (.I(\as2650.holding_reg[5] ),
    .Z(_1056_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5652_ (.I(_0917_),
    .Z(_1057_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5653_ (.A1(_1056_),
    .A2(_1057_),
    .ZN(_1058_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5654_ (.A1(_1055_),
    .A2(_4379_),
    .B(_1058_),
    .ZN(_1059_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5655_ (.A1(_4106_),
    .A2(_0587_),
    .ZN(_1060_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _5656_ (.A1(_4115_),
    .A2(_0540_),
    .B(_1060_),
    .C(_4376_),
    .ZN(_1061_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5657_ (.A1(\as2650.holding_reg[5] ),
    .A2(_0595_),
    .B(_1061_),
    .ZN(_1062_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5658_ (.A1(_4116_),
    .A2(_0840_),
    .ZN(_1063_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5659_ (.A1(_1056_),
    .A2(_0840_),
    .B(_1063_),
    .ZN(_1064_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5660_ (.A1(_1062_),
    .A2(_1064_),
    .Z(_1065_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5661_ (.I(_1065_),
    .Z(_1066_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5662_ (.A1(_0994_),
    .A2(_1002_),
    .B(_0992_),
    .ZN(_1067_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5663_ (.A1(_1066_),
    .A2(_1067_),
    .Z(_1068_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5664_ (.A1(_1056_),
    .A2(_1061_),
    .A3(_1063_),
    .ZN(_1069_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5665_ (.A1(_1062_),
    .A2(_1064_),
    .Z(_1070_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _5666_ (.A1(_0626_),
    .A2(_1069_),
    .B1(_1070_),
    .B2(_0632_),
    .C(_0582_),
    .ZN(_1071_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5667_ (.A1(_0855_),
    .A2(_1066_),
    .B(_1071_),
    .ZN(_1072_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5668_ (.A1(_0986_),
    .A2(_0991_),
    .ZN(_1073_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5669_ (.A1(_0995_),
    .A2(_0999_),
    .B(_1073_),
    .ZN(_1074_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5670_ (.A1(_1066_),
    .A2(_1074_),
    .Z(_1075_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5671_ (.A1(_0931_),
    .A2(_1075_),
    .ZN(_1076_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5672_ (.A1(_1004_),
    .A2(_1068_),
    .B(_1072_),
    .C(_1076_),
    .ZN(_1077_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5673_ (.A1(_0583_),
    .A2(_1059_),
    .B(_1077_),
    .ZN(_1078_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _5674_ (.A1(_4172_),
    .A2(_4175_),
    .A3(_4133_),
    .A4(_0942_),
    .ZN(_1079_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5675_ (.A1(_4126_),
    .A2(_1011_),
    .B(_4116_),
    .ZN(_1080_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5676_ (.A1(_1079_),
    .A2(_1080_),
    .ZN(_1081_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _5677_ (.A1(_4115_),
    .A2(_4125_),
    .A3(_0869_),
    .A4(_4199_),
    .ZN(_1082_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _5678_ (.A1(_0951_),
    .A2(_4177_),
    .A3(_4178_),
    .B(_4173_),
    .ZN(_1083_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _5679_ (.A1(_1082_),
    .A2(_1083_),
    .A3(_0892_),
    .Z(_1084_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _5680_ (.A1(_1055_),
    .A2(_1010_),
    .B1(_1081_),
    .B2(_0941_),
    .C(_1084_),
    .ZN(_1085_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5681_ (.I(_1085_),
    .Z(_1086_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5682_ (.I(_4106_),
    .Z(_1087_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5683_ (.I(_1087_),
    .Z(_1088_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5684_ (.I(_4104_),
    .Z(_1089_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5685_ (.I(_1089_),
    .Z(_1090_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5686_ (.I(net1),
    .Z(_1091_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5687_ (.I(_1091_),
    .Z(_1092_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5688_ (.I(_1092_),
    .Z(_1093_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5689_ (.I(_1093_),
    .Z(_1094_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5690_ (.I(_1094_),
    .Z(_1095_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5691_ (.A1(_4204_),
    .A2(_1024_),
    .ZN(_1096_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5692_ (.A1(_1095_),
    .A2(_0788_),
    .B(_1096_),
    .C(_1026_),
    .ZN(_1097_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5693_ (.A1(_1090_),
    .A2(_0523_),
    .B(_1097_),
    .C(_0669_),
    .ZN(_1098_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5694_ (.I(_4189_),
    .Z(_1099_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5695_ (.A1(_1099_),
    .A2(_0783_),
    .B(_0779_),
    .ZN(_1100_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5696_ (.A1(_1088_),
    .A2(_0779_),
    .B1(_1098_),
    .B2(_1100_),
    .ZN(_1101_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _5697_ (.A1(_1082_),
    .A2(_1083_),
    .A3(_0871_),
    .Z(_1102_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _5698_ (.A1(_1055_),
    .A2(_0959_),
    .B1(_1081_),
    .B2(_1032_),
    .C(_1102_),
    .ZN(_1103_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5699_ (.I(_1103_),
    .Z(_1104_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5700_ (.A1(_1016_),
    .A2(_1104_),
    .ZN(_1105_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5701_ (.A1(_1016_),
    .A2(_1101_),
    .B(_1105_),
    .C(_0644_),
    .ZN(_1106_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5702_ (.A1(_0644_),
    .A2(_1086_),
    .B(_1106_),
    .C(_0913_),
    .ZN(_1107_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5703_ (.A1(_0748_),
    .A2(_1078_),
    .B(_1107_),
    .ZN(_1108_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5704_ (.A1(\as2650.stack[1][13] ),
    .A2(_0704_),
    .B1(_0710_),
    .B2(\as2650.stack[0][13] ),
    .ZN(_1109_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5705_ (.I(_1109_),
    .ZN(_1110_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _5706_ (.A1(\as2650.stack[3][13] ),
    .A2(_0821_),
    .B1(_0718_),
    .B2(\as2650.stack[2][13] ),
    .C(_1110_),
    .ZN(_1111_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5707_ (.A1(\as2650.stack[7][13] ),
    .A2(_1043_),
    .B1(_1044_),
    .B2(\as2650.stack[6][13] ),
    .ZN(_1112_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _5708_ (.A1(\as2650.stack[5][13] ),
    .A2(_0824_),
    .B1(_0827_),
    .B2(\as2650.stack[4][13] ),
    .C(_0825_),
    .ZN(_1113_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _5709_ (.A1(_0831_),
    .A2(_1111_),
    .B1(_1112_),
    .B2(_1113_),
    .ZN(_1114_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5710_ (.A1(_0817_),
    .A2(_1114_),
    .ZN(_1115_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5711_ (.A1(_1088_),
    .A2(_0734_),
    .ZN(_1116_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5712_ (.A1(_0742_),
    .A2(_1115_),
    .A3(_1116_),
    .ZN(_1117_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5713_ (.A1(_0579_),
    .A2(_1108_),
    .B(_1117_),
    .C(_0745_),
    .ZN(_1118_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5714_ (.A1(_1054_),
    .A2(_0983_),
    .B(_1118_),
    .ZN(_0027_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5715_ (.I(\as2650.r123[0][6] ),
    .ZN(_1119_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5716_ (.I(_4100_),
    .Z(_1120_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5717_ (.I(_1120_),
    .Z(_1121_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5718_ (.I(_1121_),
    .ZN(_1122_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5719_ (.A1(_1122_),
    .A2(_0818_),
    .ZN(_1123_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5720_ (.A1(\as2650.stack[5][14] ),
    .A2(_0705_),
    .B1(_0711_),
    .B2(\as2650.stack[4][14] ),
    .ZN(_1124_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _5721_ (.A1(\as2650.stack[7][14] ),
    .A2(_1043_),
    .B1(_1044_),
    .B2(\as2650.stack[6][14] ),
    .C(_1047_),
    .ZN(_1125_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5722_ (.A1(\as2650.stack[1][14] ),
    .A2(_0705_),
    .B1(_0711_),
    .B2(\as2650.stack[0][14] ),
    .ZN(_1126_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _5723_ (.A1(\as2650.stack[3][14] ),
    .A2(_1043_),
    .B1(_1044_),
    .B2(\as2650.stack[2][14] ),
    .C(_0973_),
    .ZN(_1127_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _5724_ (.A1(_1124_),
    .A2(_1125_),
    .B1(_1126_),
    .B2(_1127_),
    .ZN(_1128_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5725_ (.A1(_0820_),
    .A2(_1128_),
    .ZN(_1129_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5726_ (.A1(_0743_),
    .A2(_1129_),
    .ZN(_1130_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5727_ (.I(_4094_),
    .Z(_1131_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _5728_ (.A1(_0523_),
    .A2(_0652_),
    .A3(_0808_),
    .A4(_0569_),
    .ZN(_1132_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5729_ (.A1(_1131_),
    .A2(_1132_),
    .ZN(_1133_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5730_ (.A1(_4185_),
    .A2(_1079_),
    .Z(_1134_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5731_ (.A1(_1082_),
    .A2(_4102_),
    .Z(_1135_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5732_ (.A1(_0799_),
    .A2(_1135_),
    .ZN(_1136_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _5733_ (.A1(_4104_),
    .A2(_0959_),
    .B1(_1134_),
    .B2(_1032_),
    .C(_1136_),
    .ZN(_1137_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5734_ (.I(_1137_),
    .Z(_1138_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5735_ (.I(_0672_),
    .Z(_1139_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5736_ (.I(net2),
    .Z(_1140_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5737_ (.I(_1140_),
    .Z(_1141_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5738_ (.I(_1141_),
    .Z(_1142_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5739_ (.I(_1142_),
    .Z(_1143_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5740_ (.A1(_4104_),
    .A2(_4187_),
    .Z(_1144_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5741_ (.A1(_1144_),
    .A2(_0683_),
    .ZN(_1145_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5742_ (.A1(_1143_),
    .A2(_1024_),
    .B(_1145_),
    .C(_0685_),
    .ZN(_1146_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5743_ (.A1(_1139_),
    .A2(_1026_),
    .B(_1146_),
    .C(_0879_),
    .ZN(_1147_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5744_ (.A1(_1028_),
    .A2(_0669_),
    .B(_1147_),
    .C(_0689_),
    .ZN(_1148_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5745_ (.A1(_1121_),
    .A2(_0664_),
    .ZN(_1149_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5746_ (.A1(_1148_),
    .A2(_1149_),
    .B(_0781_),
    .ZN(_1150_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5747_ (.A1(_0781_),
    .A2(_1138_),
    .B(_1150_),
    .C(_0899_),
    .ZN(_1151_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5748_ (.A1(_0648_),
    .A2(_1135_),
    .ZN(_1152_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _5749_ (.A1(_4181_),
    .A2(_1010_),
    .B1(_1134_),
    .B2(_0941_),
    .C(_1152_),
    .ZN(_1153_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5750_ (.I(_1153_),
    .Z(_1154_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5751_ (.A1(_0643_),
    .A2(_1154_),
    .ZN(_1155_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5752_ (.A1(_1151_),
    .A2(_1155_),
    .ZN(_1156_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5753_ (.A1(_4100_),
    .A2(_0541_),
    .ZN(_1157_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5754_ (.A1(_4103_),
    .A2(_0541_),
    .B(_1157_),
    .C(_4378_),
    .ZN(_1158_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5755_ (.A1(_4181_),
    .A2(_4396_),
    .ZN(_1159_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5756_ (.A1(\as2650.holding_reg[6] ),
    .A2(_1158_),
    .A3(_1159_),
    .ZN(_1160_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5757_ (.A1(\as2650.holding_reg[6] ),
    .A2(_1057_),
    .B(_1158_),
    .ZN(_1161_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5758_ (.A1(\as2650.holding_reg[6] ),
    .A2(_4397_),
    .B(_1159_),
    .ZN(_1162_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5759_ (.A1(_1161_),
    .A2(_1162_),
    .ZN(_1163_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5760_ (.A1(_1160_),
    .A2(_1163_),
    .ZN(_1164_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5761_ (.I(_1164_),
    .Z(_1165_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5762_ (.A1(_1062_),
    .A2(_1059_),
    .Z(_1166_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5763_ (.A1(_1066_),
    .A2(_1074_),
    .B(_1166_),
    .ZN(_1167_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5764_ (.A1(_1165_),
    .A2(_1167_),
    .B(_0930_),
    .ZN(_1168_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5765_ (.A1(_1165_),
    .A2(_1167_),
    .B(_1168_),
    .ZN(_1169_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5766_ (.A1(_1069_),
    .A2(_1067_),
    .B(_1070_),
    .ZN(_1170_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5767_ (.A1(_1165_),
    .A2(_1170_),
    .Z(_1171_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5768_ (.A1(_1004_),
    .A2(_1171_),
    .ZN(_1172_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5769_ (.A1(_1161_),
    .A2(_1162_),
    .ZN(_1173_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _5770_ (.A1(_0625_),
    .A2(_1173_),
    .B1(_1163_),
    .B2(_1005_),
    .C(_0914_),
    .ZN(_1174_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5771_ (.A1(_0770_),
    .A2(_1165_),
    .B(_1174_),
    .ZN(_1175_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5772_ (.I(_1162_),
    .ZN(_1176_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _5773_ (.A1(_1169_),
    .A2(_1172_),
    .A3(_1175_),
    .B1(_1176_),
    .B2(_0583_),
    .ZN(_1177_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5774_ (.A1(_0694_),
    .A2(_1177_),
    .ZN(_1178_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _5775_ (.A1(_0913_),
    .A2(_1156_),
    .B(_1178_),
    .ZN(_1179_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5776_ (.A1(_1133_),
    .A2(_1179_),
    .ZN(_1180_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5777_ (.A1(_1123_),
    .A2(_1130_),
    .B(_0745_),
    .C(_1180_),
    .ZN(_1181_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5778_ (.A1(_1119_),
    .A2(_0983_),
    .B(_1181_),
    .ZN(_0028_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5779_ (.I(\as2650.r123[0][7] ),
    .ZN(_1182_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5780_ (.A1(\as2650.holding_reg[7] ),
    .A2(_1057_),
    .ZN(_1183_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5781_ (.A1(_0671_),
    .A2(_1057_),
    .B(_1183_),
    .ZN(_1184_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _5782_ (.I(_1184_),
    .ZN(_1185_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5783_ (.I(_4076_),
    .Z(_1186_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5784_ (.I(_1186_),
    .Z(_1187_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5785_ (.A1(_0670_),
    .A2(_0640_),
    .ZN(_1188_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _5786_ (.A1(_1187_),
    .A2(_0640_),
    .B(_1188_),
    .C(_4379_),
    .ZN(_1189_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5787_ (.A1(\as2650.holding_reg[7] ),
    .A2(_4397_),
    .ZN(_1190_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5788_ (.A1(_1189_),
    .A2(_1190_),
    .ZN(_1191_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5789_ (.A1(_1191_),
    .A2(_1184_),
    .ZN(_1192_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5790_ (.A1(_1189_),
    .A2(_1190_),
    .A3(_1185_),
    .ZN(_1193_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5791_ (.A1(_1192_),
    .A2(_1193_),
    .ZN(_1194_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5792_ (.I(_1194_),
    .Z(_1195_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5793_ (.A1(_1173_),
    .A2(_1170_),
    .B(_1163_),
    .ZN(_1196_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5794_ (.A1(_1195_),
    .A2(_1196_),
    .B(_0616_),
    .ZN(_1197_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5795_ (.A1(_1195_),
    .A2(_1196_),
    .B(_1197_),
    .ZN(_1198_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5796_ (.A1(_1189_),
    .A2(_1190_),
    .B(_1185_),
    .ZN(_1199_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5797_ (.A1(_1191_),
    .A2(_1184_),
    .ZN(_1200_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5798_ (.A1(_1199_),
    .A2(_1200_),
    .ZN(_1201_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5799_ (.A1(_1161_),
    .A2(_1176_),
    .ZN(_1202_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5800_ (.A1(_1164_),
    .A2(_1167_),
    .B(_1202_),
    .ZN(_1203_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5801_ (.A1(_1201_),
    .A2(_1203_),
    .Z(_1204_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _5802_ (.A1(_0625_),
    .A2(_1199_),
    .B1(_1193_),
    .B2(_1005_),
    .C(_0856_),
    .ZN(_1205_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5803_ (.A1(_0628_),
    .A2(_1195_),
    .B(_1205_),
    .ZN(_1206_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5804_ (.A1(_0930_),
    .A2(_1204_),
    .B(_1206_),
    .ZN(_1207_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _5805_ (.A1(_0914_),
    .A2(_1185_),
    .B1(_1198_),
    .B2(_1207_),
    .ZN(_1208_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5806_ (.I(_1208_),
    .Z(_1209_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5807_ (.I(_1187_),
    .Z(_1210_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5808_ (.I(_1210_),
    .Z(_1211_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5809_ (.I(_0609_),
    .Z(_1212_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5810_ (.A1(_1212_),
    .A2(_0782_),
    .B(_0612_),
    .ZN(_1213_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _5811_ (.I(net3),
    .ZN(_1214_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5812_ (.I(_1214_),
    .Z(_1215_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5813_ (.I(_1215_),
    .Z(_1216_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5814_ (.I(_4184_),
    .Z(_1217_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5815_ (.A1(_1217_),
    .A2(_0682_),
    .ZN(_1218_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5816_ (.A1(_1216_),
    .A2(_1024_),
    .B(_1218_),
    .C(_0685_),
    .ZN(_1219_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5817_ (.A1(_1026_),
    .A2(_1213_),
    .B(_1219_),
    .C(_0879_),
    .ZN(_1220_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5818_ (.A1(_1089_),
    .A2(_0669_),
    .B(_1220_),
    .C(_0689_),
    .ZN(_1221_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5819_ (.A1(_1211_),
    .A2(_0878_),
    .B(_0661_),
    .C(_1221_),
    .ZN(_1222_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5820_ (.A1(_4181_),
    .A2(_1079_),
    .ZN(_1223_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5821_ (.A1(_0671_),
    .A2(_1223_),
    .Z(_1224_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5822_ (.A1(_4179_),
    .A2(_4103_),
    .ZN(_1225_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5823_ (.A1(_4081_),
    .A2(_1225_),
    .Z(_1226_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _5824_ (.A1(_0672_),
    .A2(_0959_),
    .B1(_1224_),
    .B2(_1032_),
    .C1(_1226_),
    .C2(_0871_),
    .ZN(_1227_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5825_ (.I(_1227_),
    .Z(_1228_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5826_ (.A1(_0781_),
    .A2(_1228_),
    .ZN(_1229_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5827_ (.A1(_0692_),
    .A2(_1222_),
    .A3(_1229_),
    .ZN(_1230_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5828_ (.A1(_0941_),
    .A2(_1224_),
    .ZN(_1231_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5829_ (.A1(_0671_),
    .A2(_1010_),
    .B1(_1226_),
    .B2(_0892_),
    .ZN(_1232_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5830_ (.A1(_1231_),
    .A2(_1232_),
    .ZN(_1233_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5831_ (.I(_1233_),
    .Z(_1234_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5832_ (.A1(_0899_),
    .A2(_1234_),
    .ZN(_1235_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5833_ (.A1(_1230_),
    .A2(_1235_),
    .ZN(_1236_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5834_ (.A1(_0580_),
    .A2(_1236_),
    .ZN(_1237_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5835_ (.A1(_0748_),
    .A2(_1209_),
    .B(_1237_),
    .ZN(_1238_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5836_ (.A1(_1133_),
    .A2(_1238_),
    .Z(_1239_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5837_ (.I(_1211_),
    .Z(_1240_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5838_ (.A1(_1240_),
    .A2(_0818_),
    .Z(_1241_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5839_ (.A1(_0744_),
    .A2(_1241_),
    .B(_0577_),
    .ZN(_1242_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5840_ (.A1(_1182_),
    .A2(_0983_),
    .B1(_1239_),
    .B2(_1242_),
    .ZN(_0029_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5841_ (.I(_0720_),
    .Z(_1243_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5842_ (.A1(_4238_),
    .A2(_4288_),
    .ZN(_1244_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5843_ (.I(_1244_),
    .Z(_1245_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _5844_ (.I(\as2650.cycle[0] ),
    .ZN(_1246_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5845_ (.A1(_1246_),
    .A2(_0347_),
    .ZN(_1247_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5846_ (.A1(\as2650.halted ),
    .A2(_1247_),
    .ZN(_1248_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _5847_ (.A1(_0494_),
    .A2(_0630_),
    .B(_4316_),
    .ZN(_1249_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5848_ (.A1(_4358_),
    .A2(_0390_),
    .ZN(_1250_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _5849_ (.A1(_0396_),
    .A2(_1248_),
    .A3(_1249_),
    .A4(_1250_),
    .ZN(_1251_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5850_ (.A1(_4046_),
    .A2(_1246_),
    .ZN(_1252_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5851_ (.A1(_0341_),
    .A2(_1252_),
    .ZN(_1253_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5852_ (.A1(_0460_),
    .A2(_1249_),
    .ZN(_1254_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5853_ (.A1(_0614_),
    .A2(_0359_),
    .B1(_1245_),
    .B2(_1254_),
    .ZN(_1255_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _5854_ (.A1(_4243_),
    .A2(_0462_),
    .A3(_1253_),
    .A4(_1255_),
    .ZN(_1256_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5855_ (.A1(_1245_),
    .A2(_1251_),
    .B(_1256_),
    .ZN(_1257_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5856_ (.I(_4279_),
    .Z(_1258_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5857_ (.I(_0527_),
    .Z(_1259_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5858_ (.A1(_0337_),
    .A2(_4245_),
    .A3(_1259_),
    .ZN(_1260_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5859_ (.A1(_4439_),
    .A2(_0341_),
    .A3(_0442_),
    .ZN(_1261_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _5860_ (.A1(_4285_),
    .A2(_1249_),
    .A3(_1260_),
    .A4(_1261_),
    .ZN(_1262_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5861_ (.A1(_4391_),
    .A2(_1258_),
    .B(_1262_),
    .ZN(_1263_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5862_ (.I(_0474_),
    .Z(_1264_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5863_ (.A1(_1131_),
    .A2(_0367_),
    .A3(_1264_),
    .ZN(_1265_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5864_ (.A1(_4358_),
    .A2(_0556_),
    .ZN(_1266_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _5865_ (.A1(_4246_),
    .A2(_1265_),
    .A3(_1266_),
    .ZN(_1267_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _5866_ (.A1(_4343_),
    .A2(_1257_),
    .B(_1263_),
    .C(_1267_),
    .ZN(_1268_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5867_ (.I(_1268_),
    .ZN(_1269_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5868_ (.I(_1269_),
    .Z(_1270_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5869_ (.A1(_1243_),
    .A2(_0719_),
    .A3(_1270_),
    .ZN(_1271_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5870_ (.I(_1271_),
    .Z(_1272_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5871_ (.I(_1267_),
    .Z(_1273_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5872_ (.I(\as2650.pc[0] ),
    .Z(_1274_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5873_ (.I(_1274_),
    .Z(_1275_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5874_ (.I(_1275_),
    .Z(_1276_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5875_ (.I(_1276_),
    .Z(_1277_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5876_ (.A1(_4045_),
    .A2(_1247_),
    .ZN(_1278_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5877_ (.I(_1278_),
    .Z(_1279_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5878_ (.A1(_4364_),
    .A2(_0479_),
    .A3(_1279_),
    .ZN(_1280_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5879_ (.I(_1280_),
    .Z(_1281_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5880_ (.A1(_1277_),
    .A2(_1281_),
    .Z(_1282_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5881_ (.A1(_0698_),
    .A2(_1273_),
    .B(_1282_),
    .ZN(_1283_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5882_ (.I(_1283_),
    .Z(_1284_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5883_ (.I(_1271_),
    .Z(_1285_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5884_ (.A1(\as2650.stack[3][0] ),
    .A2(_1285_),
    .ZN(_1286_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5885_ (.A1(_1272_),
    .A2(_1284_),
    .B(_1286_),
    .ZN(_0030_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _5886_ (.I(\as2650.pc[1] ),
    .ZN(_1287_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5887_ (.I(_1287_),
    .Z(_1288_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5888_ (.I0(_0753_),
    .I1(_1288_),
    .S(_1281_),
    .Z(_1289_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5889_ (.I(_1289_),
    .Z(_1290_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5890_ (.A1(\as2650.stack[3][1] ),
    .A2(_1285_),
    .ZN(_1291_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5891_ (.A1(_1272_),
    .A2(_1290_),
    .B(_1291_),
    .ZN(_0031_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _5892_ (.I(\as2650.pc[2] ),
    .ZN(_1292_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5893_ (.I0(_0845_),
    .I1(_1292_),
    .S(_1281_),
    .Z(_1293_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5894_ (.I(_1293_),
    .Z(_1294_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5895_ (.A1(\as2650.stack[3][2] ),
    .A2(_1285_),
    .ZN(_1295_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5896_ (.A1(_1272_),
    .A2(_1294_),
    .B(_1295_),
    .ZN(_0032_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _5897_ (.I(\as2650.pc[3] ),
    .ZN(_1296_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5898_ (.I(_1296_),
    .Z(_1297_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5899_ (.I(_1297_),
    .Z(_1298_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5900_ (.I0(_0970_),
    .I1(_1298_),
    .S(_1281_),
    .Z(_1299_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5901_ (.I(_1299_),
    .Z(_1300_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5902_ (.A1(\as2650.stack[3][3] ),
    .A2(_1285_),
    .ZN(_1301_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5903_ (.A1(_1272_),
    .A2(_1300_),
    .B(_1301_),
    .ZN(_0033_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5904_ (.I(_1271_),
    .Z(_1302_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5905_ (.I(_1018_),
    .Z(_1303_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _5906_ (.I(\as2650.pc[4] ),
    .ZN(_1304_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5907_ (.I(_1304_),
    .Z(_1305_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5908_ (.I(_1267_),
    .Z(_1306_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5909_ (.A1(_1305_),
    .A2(_1306_),
    .ZN(_1307_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5910_ (.A1(_1303_),
    .A2(_1273_),
    .B(_1307_),
    .ZN(_1308_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5911_ (.I(_1308_),
    .Z(_1309_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5912_ (.I(_1271_),
    .Z(_1310_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5913_ (.A1(\as2650.stack[3][4] ),
    .A2(_1310_),
    .ZN(_1311_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5914_ (.A1(_1302_),
    .A2(_1309_),
    .B(_1311_),
    .ZN(_0034_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5915_ (.I(_1088_),
    .Z(_1312_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _5916_ (.I(\as2650.pc[5] ),
    .ZN(_1313_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5917_ (.I(_1313_),
    .Z(_1314_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5918_ (.A1(_1314_),
    .A2(_1306_),
    .ZN(_1315_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5919_ (.A1(_1312_),
    .A2(_1273_),
    .B(_1315_),
    .ZN(_1316_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5920_ (.I(_1316_),
    .Z(_1317_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5921_ (.A1(\as2650.stack[3][5] ),
    .A2(_1310_),
    .ZN(_1318_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5922_ (.A1(_1302_),
    .A2(_1317_),
    .B(_1318_),
    .ZN(_0035_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5923_ (.I(_1121_),
    .Z(_1319_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5924_ (.I(\as2650.pc[6] ),
    .Z(_1320_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5925_ (.I(_1320_),
    .Z(_1321_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5926_ (.I(_1321_),
    .Z(_1322_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5927_ (.A1(_1322_),
    .A2(_1280_),
    .Z(_1323_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5928_ (.A1(_1319_),
    .A2(_1273_),
    .B(_1323_),
    .ZN(_1324_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5929_ (.I(_1324_),
    .Z(_1325_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5930_ (.A1(\as2650.stack[3][6] ),
    .A2(_1310_),
    .ZN(_1326_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5931_ (.A1(_1302_),
    .A2(_1325_),
    .B(_1326_),
    .ZN(_0036_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _5932_ (.I(\as2650.pc[7] ),
    .ZN(_1327_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5933_ (.I(_1327_),
    .Z(_1328_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5934_ (.A1(_1328_),
    .A2(_1306_),
    .ZN(_1329_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5935_ (.A1(_1211_),
    .A2(_1306_),
    .B(_1329_),
    .ZN(_1330_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5936_ (.I(_1330_),
    .Z(_1331_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5937_ (.A1(\as2650.stack[3][7] ),
    .A2(_1310_),
    .ZN(_1332_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5938_ (.A1(_1302_),
    .A2(_1331_),
    .B(_1332_),
    .ZN(_0037_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5939_ (.A1(_1243_),
    .A2(_0705_),
    .A3(_1270_),
    .ZN(_1333_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5940_ (.I(_1333_),
    .Z(_1334_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5941_ (.I(_1333_),
    .Z(_1335_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5942_ (.A1(\as2650.stack[2][0] ),
    .A2(_1335_),
    .ZN(_1336_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5943_ (.A1(_1284_),
    .A2(_1334_),
    .B(_1336_),
    .ZN(_0038_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5944_ (.A1(\as2650.stack[2][1] ),
    .A2(_1335_),
    .ZN(_1337_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5945_ (.A1(_1290_),
    .A2(_1334_),
    .B(_1337_),
    .ZN(_0039_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5946_ (.A1(\as2650.stack[2][2] ),
    .A2(_1335_),
    .ZN(_1338_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5947_ (.A1(_1294_),
    .A2(_1334_),
    .B(_1338_),
    .ZN(_0040_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5948_ (.A1(\as2650.stack[2][3] ),
    .A2(_1335_),
    .ZN(_1339_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5949_ (.A1(_1300_),
    .A2(_1334_),
    .B(_1339_),
    .ZN(_0041_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5950_ (.I(_1333_),
    .Z(_1340_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5951_ (.I(_1333_),
    .Z(_1341_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5952_ (.A1(\as2650.stack[2][4] ),
    .A2(_1341_),
    .ZN(_1342_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5953_ (.A1(_1309_),
    .A2(_1340_),
    .B(_1342_),
    .ZN(_0042_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5954_ (.A1(\as2650.stack[2][5] ),
    .A2(_1341_),
    .ZN(_1343_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5955_ (.A1(_1317_),
    .A2(_1340_),
    .B(_1343_),
    .ZN(_0043_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5956_ (.A1(\as2650.stack[2][6] ),
    .A2(_1341_),
    .ZN(_1344_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5957_ (.A1(_1325_),
    .A2(_1340_),
    .B(_1344_),
    .ZN(_0044_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5958_ (.A1(\as2650.stack[2][7] ),
    .A2(_1341_),
    .ZN(_1345_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5959_ (.A1(_1331_),
    .A2(_1340_),
    .B(_1345_),
    .ZN(_0045_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5960_ (.I(_0700_),
    .Z(_1346_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5961_ (.I(_1269_),
    .Z(_1347_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5962_ (.I(_0708_),
    .Z(_1348_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5963_ (.I(_1348_),
    .Z(_1349_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5964_ (.I(\as2650.psu[2] ),
    .Z(_1350_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5965_ (.I(_1350_),
    .Z(_1351_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5966_ (.A1(_1349_),
    .A2(_1351_),
    .ZN(_1352_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5967_ (.A1(_1346_),
    .A2(_1347_),
    .A3(_1352_),
    .ZN(_1353_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5968_ (.I(_1353_),
    .Z(_1354_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5969_ (.I(_1353_),
    .Z(_1355_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5970_ (.A1(\as2650.stack[1][0] ),
    .A2(_1355_),
    .ZN(_1356_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5971_ (.A1(_1284_),
    .A2(_1354_),
    .B(_1356_),
    .ZN(_0046_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5972_ (.A1(\as2650.stack[1][1] ),
    .A2(_1355_),
    .ZN(_1357_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5973_ (.A1(_1290_),
    .A2(_1354_),
    .B(_1357_),
    .ZN(_0047_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5974_ (.A1(\as2650.stack[1][2] ),
    .A2(_1355_),
    .ZN(_1358_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5975_ (.A1(_1294_),
    .A2(_1354_),
    .B(_1358_),
    .ZN(_0048_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5976_ (.A1(\as2650.stack[1][3] ),
    .A2(_1355_),
    .ZN(_1359_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5977_ (.A1(_1300_),
    .A2(_1354_),
    .B(_1359_),
    .ZN(_0049_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5978_ (.I(_1353_),
    .Z(_1360_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5979_ (.I(_1353_),
    .Z(_1361_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5980_ (.A1(\as2650.stack[1][4] ),
    .A2(_1361_),
    .ZN(_1362_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5981_ (.A1(_1309_),
    .A2(_1360_),
    .B(_1362_),
    .ZN(_0050_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5982_ (.A1(\as2650.stack[1][5] ),
    .A2(_1361_),
    .ZN(_1363_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5983_ (.A1(_1317_),
    .A2(_1360_),
    .B(_1363_),
    .ZN(_0051_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5984_ (.A1(\as2650.stack[1][6] ),
    .A2(_1361_),
    .ZN(_1364_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5985_ (.A1(_1325_),
    .A2(_1360_),
    .B(_1364_),
    .ZN(_0052_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5986_ (.A1(\as2650.stack[1][7] ),
    .A2(_1361_),
    .ZN(_1365_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5987_ (.A1(_1331_),
    .A2(_1360_),
    .B(_1365_),
    .ZN(_0053_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5988_ (.I(_1350_),
    .Z(_1366_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5989_ (.I(_1268_),
    .Z(_1367_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _5990_ (.A1(_0707_),
    .A2(_1348_),
    .A3(_1366_),
    .A4(_1367_),
    .ZN(_1368_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5991_ (.I(_1368_),
    .Z(_1369_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5992_ (.I(_1369_),
    .Z(_1370_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5993_ (.A1(_4360_),
    .A2(_0479_),
    .A3(_0560_),
    .ZN(_1371_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5994_ (.I(_1371_),
    .Z(_1372_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5995_ (.I(_1372_),
    .Z(_1373_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5996_ (.I(_1372_),
    .Z(_1374_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5997_ (.A1(_0549_),
    .A2(_1280_),
    .ZN(_1375_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5998_ (.I(_1375_),
    .Z(_1376_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5999_ (.A1(\as2650.r123_2[0][0] ),
    .A2(_1376_),
    .ZN(_1377_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6000_ (.I(\as2650.pc[8] ),
    .Z(_1378_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6001_ (.I(_1378_),
    .Z(_1379_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6002_ (.I(_1379_),
    .Z(_1380_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6003_ (.I(_1380_),
    .Z(_1381_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6004_ (.A1(_0555_),
    .A2(_1267_),
    .ZN(_1382_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6005_ (.A1(_1381_),
    .A2(_1382_),
    .ZN(_1383_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6006_ (.A1(_1374_),
    .A2(_1377_),
    .A3(_1383_),
    .ZN(_1384_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6007_ (.A1(\as2650.r123[0][0] ),
    .A2(_1373_),
    .B(_1384_),
    .ZN(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6008_ (.I(_1385_),
    .Z(_1386_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6009_ (.I(_1369_),
    .Z(_1387_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6010_ (.A1(\as2650.stack[1][8] ),
    .A2(_1387_),
    .ZN(_1388_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6011_ (.A1(_1370_),
    .A2(_1386_),
    .B(_1388_),
    .ZN(_0054_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6012_ (.I(\as2650.pc[9] ),
    .ZN(_1389_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6013_ (.I(_1389_),
    .Z(_1390_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6014_ (.I(_1375_),
    .Z(_1391_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6015_ (.I(_1371_),
    .Z(_1392_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6016_ (.A1(\as2650.r123_2[0][1] ),
    .A2(_1376_),
    .ZN(_1393_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6017_ (.A1(_1390_),
    .A2(_1391_),
    .B(_1392_),
    .C(_1393_),
    .ZN(_1394_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6018_ (.A1(\as2650.r123[0][1] ),
    .A2(_1373_),
    .B(_1394_),
    .ZN(_1395_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6019_ (.I(_1395_),
    .Z(_1396_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6020_ (.I(_1368_),
    .Z(_1397_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6021_ (.A1(\as2650.stack[1][9] ),
    .A2(_1397_),
    .ZN(_1398_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6022_ (.A1(_1370_),
    .A2(_1396_),
    .B(_1398_),
    .ZN(_0055_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6023_ (.I(\as2650.pc[10] ),
    .ZN(_1399_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6024_ (.I(_1399_),
    .Z(_1400_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6025_ (.A1(\as2650.r123_2[0][2] ),
    .A2(_1375_),
    .ZN(_1401_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6026_ (.A1(_1400_),
    .A2(_1391_),
    .B(_1372_),
    .C(_1401_),
    .ZN(_1402_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6027_ (.A1(\as2650.r123[0][2] ),
    .A2(_1373_),
    .B(_1402_),
    .ZN(_1403_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6028_ (.I(_1403_),
    .Z(_1404_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6029_ (.A1(\as2650.stack[1][10] ),
    .A2(_1397_),
    .ZN(_1405_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6030_ (.A1(_1370_),
    .A2(_1404_),
    .B(_1405_),
    .ZN(_0056_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6031_ (.I(\as2650.pc[11] ),
    .Z(_1406_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6032_ (.I(_1406_),
    .Z(_1407_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6033_ (.I(_1407_),
    .Z(_1408_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6034_ (.I(_1408_),
    .Z(_1409_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6035_ (.A1(_1409_),
    .A2(_1382_),
    .ZN(_1410_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6036_ (.A1(\as2650.r123_2[0][3] ),
    .A2(_1391_),
    .ZN(_1411_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6037_ (.A1(_1392_),
    .A2(_1410_),
    .A3(_1411_),
    .ZN(_1412_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6038_ (.A1(\as2650.r123[0][3] ),
    .A2(_1373_),
    .B(_1412_),
    .ZN(_1413_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6039_ (.I(_1413_),
    .Z(_1414_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6040_ (.A1(\as2650.stack[1][11] ),
    .A2(_1397_),
    .ZN(_1415_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6041_ (.A1(_1370_),
    .A2(_1414_),
    .B(_1415_),
    .ZN(_0057_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _6042_ (.I(\as2650.pc[12] ),
    .ZN(_1416_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6043_ (.A1(\as2650.r123_2[0][4] ),
    .A2(_1375_),
    .ZN(_1417_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6044_ (.A1(_1416_),
    .A2(_1391_),
    .B(_1372_),
    .C(_1417_),
    .ZN(_1418_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6045_ (.A1(\as2650.r123[0][4] ),
    .A2(_1374_),
    .B(_1418_),
    .ZN(_1419_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6046_ (.I(_1419_),
    .Z(_1420_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6047_ (.A1(\as2650.stack[1][12] ),
    .A2(_1397_),
    .ZN(_1421_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6048_ (.A1(_1387_),
    .A2(_1420_),
    .B(_1421_),
    .ZN(_0058_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6049_ (.I(\as2650.pc[13] ),
    .Z(_1422_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6050_ (.A1(_1422_),
    .A2(_1382_),
    .ZN(_1423_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6051_ (.A1(\as2650.r123_2[0][5] ),
    .A2(_1376_),
    .ZN(_1424_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6052_ (.A1(_1392_),
    .A2(_1423_),
    .A3(_1424_),
    .ZN(_1425_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6053_ (.A1(\as2650.r123[0][5] ),
    .A2(_1374_),
    .B(_1425_),
    .ZN(_1426_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6054_ (.I(_1426_),
    .Z(_1427_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6055_ (.A1(\as2650.stack[1][13] ),
    .A2(_1369_),
    .ZN(_1428_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6056_ (.A1(_1387_),
    .A2(_1427_),
    .B(_1428_),
    .ZN(_0059_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6057_ (.I(\as2650.pc[14] ),
    .Z(_1429_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6058_ (.A1(_1429_),
    .A2(_1382_),
    .ZN(_1430_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6059_ (.A1(\as2650.r123_2[0][6] ),
    .A2(_1376_),
    .ZN(_1431_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6060_ (.A1(_1392_),
    .A2(_1430_),
    .A3(_1431_),
    .ZN(_1432_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6061_ (.A1(\as2650.r123[0][6] ),
    .A2(_1374_),
    .B(_1432_),
    .ZN(_1433_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6062_ (.I(_1433_),
    .Z(_1434_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6063_ (.A1(\as2650.stack[1][14] ),
    .A2(_1369_),
    .ZN(_1435_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6064_ (.A1(_1387_),
    .A2(_1434_),
    .B(_1435_),
    .ZN(_0060_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6065_ (.I(_0707_),
    .Z(_1436_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6066_ (.A1(_1436_),
    .A2(_1347_),
    .A3(_1352_),
    .ZN(_1437_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6067_ (.I(_1437_),
    .Z(_1438_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6068_ (.I(_1437_),
    .Z(_1439_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6069_ (.A1(\as2650.stack[0][0] ),
    .A2(_1439_),
    .ZN(_1440_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6070_ (.A1(_1284_),
    .A2(_1438_),
    .B(_1440_),
    .ZN(_0061_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6071_ (.A1(\as2650.stack[0][1] ),
    .A2(_1439_),
    .ZN(_1441_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6072_ (.A1(_1290_),
    .A2(_1438_),
    .B(_1441_),
    .ZN(_0062_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6073_ (.A1(\as2650.stack[0][2] ),
    .A2(_1439_),
    .ZN(_1442_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6074_ (.A1(_1294_),
    .A2(_1438_),
    .B(_1442_),
    .ZN(_0063_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6075_ (.A1(\as2650.stack[0][3] ),
    .A2(_1439_),
    .ZN(_1443_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6076_ (.A1(_1300_),
    .A2(_1438_),
    .B(_1443_),
    .ZN(_0064_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6077_ (.I(_1437_),
    .Z(_1444_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6078_ (.I(_1437_),
    .Z(_1445_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6079_ (.A1(\as2650.stack[0][4] ),
    .A2(_1445_),
    .ZN(_1446_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6080_ (.A1(_1309_),
    .A2(_1444_),
    .B(_1446_),
    .ZN(_0065_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6081_ (.A1(\as2650.stack[0][5] ),
    .A2(_1445_),
    .ZN(_1447_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6082_ (.A1(_1317_),
    .A2(_1444_),
    .B(_1447_),
    .ZN(_0066_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6083_ (.A1(\as2650.stack[0][6] ),
    .A2(_1445_),
    .ZN(_1448_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6084_ (.A1(_1325_),
    .A2(_1444_),
    .B(_1448_),
    .ZN(_0067_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6085_ (.A1(\as2650.stack[0][7] ),
    .A2(_1445_),
    .ZN(_1449_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6086_ (.A1(_1331_),
    .A2(_1444_),
    .B(_1449_),
    .ZN(_0068_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6087_ (.I(\as2650.r123_2[3][0] ),
    .Z(_1450_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6088_ (.I(_1450_),
    .Z(_0069_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6089_ (.I(\as2650.r123_2[3][1] ),
    .Z(_1451_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6090_ (.I(_1451_),
    .Z(_0070_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6091_ (.I(\as2650.r123_2[3][2] ),
    .Z(_1452_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6092_ (.I(_1452_),
    .Z(_0071_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6093_ (.I(\as2650.r123_2[3][3] ),
    .Z(_1453_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6094_ (.I(_1453_),
    .Z(_0072_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6095_ (.I(\as2650.r123_2[3][4] ),
    .Z(_1454_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6096_ (.I(_1454_),
    .Z(_0073_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6097_ (.I(\as2650.r123_2[3][5] ),
    .Z(_1455_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6098_ (.I(_1455_),
    .Z(_0074_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6099_ (.I(\as2650.r123_2[3][6] ),
    .Z(_1456_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6100_ (.I(_1456_),
    .Z(_0075_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6101_ (.I(\as2650.r123_2[3][7] ),
    .Z(_1457_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6102_ (.I(_1457_),
    .Z(_0076_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6103_ (.I(\as2650.psu[5] ),
    .ZN(_1458_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6104_ (.I(_0562_),
    .Z(_1459_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6105_ (.A1(_0731_),
    .A2(_0501_),
    .ZN(_1460_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _6106_ (.A1(_4047_),
    .A2(_0738_),
    .A3(_0485_),
    .A4(_1460_),
    .ZN(_1461_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6107_ (.A1(_1459_),
    .A2(_1461_),
    .B(_4329_),
    .ZN(_1462_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6108_ (.I(_0814_),
    .Z(_1463_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6109_ (.A1(_1463_),
    .A2(_0369_),
    .A3(_1264_),
    .ZN(_1464_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6110_ (.I(_4060_),
    .Z(_1465_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6111_ (.A1(_1465_),
    .A2(_0472_),
    .ZN(_1466_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6112_ (.A1(_4253_),
    .A2(_4295_),
    .ZN(_1467_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6113_ (.I(_4316_),
    .Z(_1468_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _6114_ (.A1(_1467_),
    .A2(_1468_),
    .A3(_0495_),
    .ZN(_1469_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6115_ (.A1(_1466_),
    .A2(_1469_),
    .B(_0736_),
    .ZN(_1470_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6116_ (.A1(_0446_),
    .A2(_1470_),
    .Z(_1471_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6117_ (.I(_0572_),
    .Z(_1472_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6118_ (.I(_0737_),
    .Z(_1473_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6119_ (.I(_1473_),
    .Z(_1474_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6120_ (.A1(_0739_),
    .A2(_1472_),
    .B(_1474_),
    .ZN(_1475_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6121_ (.A1(_1131_),
    .A2(_1469_),
    .ZN(_1476_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6122_ (.I(_0445_),
    .Z(_1477_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6123_ (.I(_0812_),
    .Z(_1478_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6124_ (.I(_1478_),
    .Z(_1479_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6125_ (.A1(_1479_),
    .A2(_0855_),
    .ZN(_1480_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6126_ (.I(_0550_),
    .Z(_1481_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6127_ (.I(_1481_),
    .Z(_1482_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _6128_ (.A1(_4243_),
    .A2(_4445_),
    .A3(_0449_),
    .A4(_1482_),
    .ZN(_1483_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6129_ (.A1(_0437_),
    .A2(_4235_),
    .B1(_1477_),
    .B2(_1480_),
    .C(_1483_),
    .ZN(_1484_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6130_ (.A1(_1475_),
    .A2(_1476_),
    .A3(_1484_),
    .ZN(_1485_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6131_ (.A1(_1471_),
    .A2(_1485_),
    .ZN(_1486_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6132_ (.A1(_1462_),
    .A2(_1464_),
    .A3(_1486_),
    .ZN(_1487_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6133_ (.I(_1478_),
    .Z(_1488_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6134_ (.I(_1488_),
    .Z(_1489_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6135_ (.I(_1095_),
    .Z(_1490_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6136_ (.A1(_1489_),
    .A2(_1490_),
    .ZN(_1491_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6137_ (.A1(_1088_),
    .A2(_4361_),
    .ZN(_1492_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6138_ (.I(_4374_),
    .Z(_1493_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _6139_ (.A1(_4298_),
    .A2(_4390_),
    .A3(_4369_),
    .A4(_0631_),
    .ZN(_1494_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6140_ (.I(_1494_),
    .Z(_1495_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6141_ (.A1(_1493_),
    .A2(_1495_),
    .ZN(_1496_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6142_ (.I(_1496_),
    .Z(_1497_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6143_ (.A1(_1492_),
    .A2(_1497_),
    .ZN(_1498_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6144_ (.I(_1488_),
    .Z(_1499_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _6145_ (.I(net1),
    .ZN(_1500_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6146_ (.I(_1500_),
    .Z(_1501_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6147_ (.I(_1501_),
    .Z(_1502_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6148_ (.A1(_1499_),
    .A2(_1502_),
    .B(_1492_),
    .ZN(_1503_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6149_ (.A1(\as2650.psu[5] ),
    .A2(_1491_),
    .B1(_1498_),
    .B2(_1503_),
    .ZN(_1504_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6150_ (.A1(_1477_),
    .A2(_1504_),
    .ZN(_1505_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6151_ (.A1(_1487_),
    .A2(_1505_),
    .ZN(_1506_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6152_ (.I(_0468_),
    .Z(_1507_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6153_ (.I(_1507_),
    .Z(_1508_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6154_ (.A1(_1458_),
    .A2(_1487_),
    .B(_1506_),
    .C(_1508_),
    .ZN(_0077_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6155_ (.I(_4342_),
    .Z(_1509_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6156_ (.I(_4300_),
    .Z(_1510_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6157_ (.A1(_4440_),
    .A2(_1510_),
    .ZN(_1511_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6158_ (.A1(_4439_),
    .A2(_0445_),
    .ZN(_1512_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6159_ (.A1(_4357_),
    .A2(_4297_),
    .ZN(_1513_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6160_ (.A1(_4345_),
    .A2(_1513_),
    .ZN(_1514_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _6161_ (.A1(_4241_),
    .A2(_1512_),
    .A3(_1248_),
    .A4(_1514_),
    .ZN(_1515_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6162_ (.A1(_4320_),
    .A2(_0364_),
    .A3(_1515_),
    .ZN(_1516_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _6163_ (.A1(_1509_),
    .A2(_4317_),
    .A3(_1511_),
    .B(_1516_),
    .ZN(_1517_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6164_ (.A1(_0383_),
    .A2(_4348_),
    .ZN(_1518_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6165_ (.A1(_4433_),
    .A2(_4344_),
    .ZN(_1519_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6166_ (.A1(_1513_),
    .A2(_1519_),
    .Z(_1520_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6167_ (.A1(_1518_),
    .A2(_1520_),
    .ZN(_1521_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6168_ (.A1(_4416_),
    .A2(_0315_),
    .Z(_1522_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _6169_ (.A1(_0385_),
    .A2(_4420_),
    .B1(_1521_),
    .B2(_1522_),
    .ZN(_1523_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6170_ (.I(_4359_),
    .Z(_1524_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6171_ (.A1(_1524_),
    .A2(_4445_),
    .A3(_0381_),
    .ZN(_1525_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6172_ (.A1(_1521_),
    .A2(_1525_),
    .Z(_1526_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6173_ (.A1(_4430_),
    .A2(_0325_),
    .B(_4335_),
    .ZN(_1527_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _6174_ (.A1(_0317_),
    .A2(_4338_),
    .B(_1521_),
    .C(_1527_),
    .ZN(_1528_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _6175_ (.A1(_1517_),
    .A2(_1523_),
    .A3(_1526_),
    .A4(_1528_),
    .ZN(_1529_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6176_ (.I(_1529_),
    .Z(_1530_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6177_ (.I(_0534_),
    .Z(_1531_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6178_ (.A1(_0385_),
    .A2(_1531_),
    .Z(_1532_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6179_ (.I(_1532_),
    .Z(_1533_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6180_ (.I(_0782_),
    .Z(_1534_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6181_ (.I(_1532_),
    .Z(_1535_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6182_ (.A1(_1534_),
    .A2(_1535_),
    .ZN(_1536_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6183_ (.A1(_0698_),
    .A2(_1533_),
    .B(_1536_),
    .ZN(_1537_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6184_ (.I(_1529_),
    .Z(_1538_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6185_ (.A1(net42),
    .A2(_1538_),
    .ZN(_1539_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6186_ (.A1(_1530_),
    .A2(_1537_),
    .B(_1539_),
    .C(_1508_),
    .ZN(_0078_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6187_ (.I(_0778_),
    .Z(_1540_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6188_ (.I(_0674_),
    .Z(_1541_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6189_ (.A1(_1541_),
    .A2(_1535_),
    .ZN(_1542_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6190_ (.A1(_1540_),
    .A2(_1533_),
    .B(_1542_),
    .ZN(_1543_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6191_ (.A1(net43),
    .A2(_1538_),
    .ZN(_1544_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6192_ (.A1(_1530_),
    .A2(_1543_),
    .B(_1544_),
    .C(_1508_),
    .ZN(_0079_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6193_ (.I(_0877_),
    .Z(_1545_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6194_ (.A1(_0950_),
    .A2(_1535_),
    .ZN(_1546_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6195_ (.A1(_1545_),
    .A2(_1533_),
    .B(_1546_),
    .ZN(_1547_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6196_ (.A1(net44),
    .A2(_1538_),
    .ZN(_1548_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6197_ (.I(_0469_),
    .Z(_1549_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6198_ (.A1(_1530_),
    .A2(_1547_),
    .B(_1548_),
    .C(_1549_),
    .ZN(_0080_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6199_ (.I(_0880_),
    .Z(_1550_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6200_ (.A1(_1550_),
    .A2(_1535_),
    .ZN(_1551_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6201_ (.A1(_0969_),
    .A2(_1533_),
    .B(_1551_),
    .ZN(_1552_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6202_ (.A1(net45),
    .A2(_1538_),
    .ZN(_1553_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6203_ (.A1(_1530_),
    .A2(_1552_),
    .B(_1553_),
    .C(_1549_),
    .ZN(_0081_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6204_ (.I(_1529_),
    .Z(_1554_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6205_ (.I(_1532_),
    .Z(_1555_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6206_ (.I(_1532_),
    .Z(_1556_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6207_ (.A1(_1099_),
    .A2(_1556_),
    .ZN(_1557_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6208_ (.A1(_1303_),
    .A2(_1555_),
    .B(_1557_),
    .ZN(_1558_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6209_ (.I(_1529_),
    .Z(_1559_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6210_ (.A1(net46),
    .A2(_1559_),
    .ZN(_1560_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6211_ (.A1(_1554_),
    .A2(_1558_),
    .B(_1560_),
    .C(_1549_),
    .ZN(_0082_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6212_ (.I(_1055_),
    .Z(_1561_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6213_ (.A1(_1561_),
    .A2(_1556_),
    .ZN(_1562_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6214_ (.A1(_1312_),
    .A2(_1555_),
    .B(_1562_),
    .ZN(_1563_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6215_ (.A1(net20),
    .A2(_1559_),
    .ZN(_1564_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6216_ (.A1(_1554_),
    .A2(_1563_),
    .B(_1564_),
    .C(_1549_),
    .ZN(_0083_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6217_ (.A1(_1090_),
    .A2(_1556_),
    .ZN(_1565_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6218_ (.A1(_1319_),
    .A2(_1555_),
    .B(_1565_),
    .ZN(_1566_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6219_ (.A1(net21),
    .A2(_1559_),
    .ZN(_1567_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6220_ (.I(_1507_),
    .Z(_1568_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6221_ (.A1(_1554_),
    .A2(_1566_),
    .B(_1567_),
    .C(_1568_),
    .ZN(_0084_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6222_ (.A1(_1139_),
    .A2(_1556_),
    .ZN(_1569_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6223_ (.A1(_1240_),
    .A2(_1555_),
    .B(_1569_),
    .ZN(_1570_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6224_ (.A1(net22),
    .A2(_1559_),
    .ZN(_1571_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6225_ (.A1(_1554_),
    .A2(_1570_),
    .B(_1571_),
    .C(_1568_),
    .ZN(_0085_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6226_ (.A1(_0699_),
    .A2(_0708_),
    .ZN(_1572_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6227_ (.I(_1572_),
    .Z(_1573_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6228_ (.I(_1573_),
    .Z(_1574_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6229_ (.A1(_1351_),
    .A2(_1574_),
    .A3(_1367_),
    .ZN(_1575_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6230_ (.I(_1575_),
    .Z(_1576_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6231_ (.I(_1576_),
    .Z(_1577_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6232_ (.I(_1576_),
    .Z(_1578_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6233_ (.A1(\as2650.stack[3][8] ),
    .A2(_1578_),
    .ZN(_1579_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6234_ (.A1(_1577_),
    .A2(_1386_),
    .B(_1579_),
    .ZN(_0086_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6235_ (.I(_1575_),
    .Z(_1580_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6236_ (.A1(\as2650.stack[3][9] ),
    .A2(_1580_),
    .ZN(_1581_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6237_ (.A1(_1577_),
    .A2(_1396_),
    .B(_1581_),
    .ZN(_0087_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6238_ (.A1(\as2650.stack[3][10] ),
    .A2(_1580_),
    .ZN(_1582_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6239_ (.A1(_1577_),
    .A2(_1404_),
    .B(_1582_),
    .ZN(_0088_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6240_ (.A1(\as2650.stack[3][11] ),
    .A2(_1580_),
    .ZN(_1583_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6241_ (.A1(_1577_),
    .A2(_1414_),
    .B(_1583_),
    .ZN(_0089_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6242_ (.A1(\as2650.stack[3][12] ),
    .A2(_1580_),
    .ZN(_1584_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6243_ (.A1(_1578_),
    .A2(_1420_),
    .B(_1584_),
    .ZN(_0090_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6244_ (.A1(\as2650.stack[3][13] ),
    .A2(_1576_),
    .ZN(_1585_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6245_ (.A1(_1578_),
    .A2(_1427_),
    .B(_1585_),
    .ZN(_0091_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6246_ (.A1(\as2650.stack[3][14] ),
    .A2(_1576_),
    .ZN(_1586_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6247_ (.A1(_1578_),
    .A2(_1434_),
    .B(_1586_),
    .ZN(_0092_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6248_ (.I(_1513_),
    .Z(_1587_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6249_ (.I(_1587_),
    .Z(_1588_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6250_ (.I(_1588_),
    .Z(_1589_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _6251_ (.A1(_0615_),
    .A2(_4392_),
    .A3(_4450_),
    .ZN(_1590_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6252_ (.A1(_0839_),
    .A2(_0865_),
    .Z(_1591_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6253_ (.A1(_0775_),
    .A2(_1591_),
    .ZN(_1592_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6254_ (.A1(_0638_),
    .A2(_0940_),
    .A3(_1592_),
    .ZN(_1593_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _6255_ (.A1(_1009_),
    .A2(_1078_),
    .A3(_1177_),
    .A4(_1593_),
    .Z(_1594_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6256_ (.A1(_1160_),
    .A2(_1163_),
    .B(_1065_),
    .ZN(_1595_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6257_ (.A1(_0995_),
    .A2(_1194_),
    .A3(_1595_),
    .ZN(_1596_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6258_ (.A1(_0606_),
    .A2(_0757_),
    .ZN(_1597_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6259_ (.A1(_0848_),
    .A2(_0853_),
    .ZN(_1598_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6260_ (.A1(_0861_),
    .A2(_1597_),
    .B(_1598_),
    .ZN(_1599_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6261_ (.A1(_0922_),
    .A2(_0923_),
    .ZN(_1600_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6262_ (.A1(_0933_),
    .A2(_1599_),
    .B(_1600_),
    .ZN(_1601_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6263_ (.A1(_0998_),
    .A2(_1601_),
    .Z(_1602_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6264_ (.A1(_1062_),
    .A2(_1059_),
    .ZN(_1603_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6265_ (.A1(_1164_),
    .A2(_1603_),
    .B1(_1595_),
    .B2(_1073_),
    .C(_1202_),
    .ZN(_1604_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6266_ (.A1(_1201_),
    .A2(_1604_),
    .ZN(_1605_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6267_ (.A1(_1191_),
    .A2(_1185_),
    .B(_1605_),
    .ZN(_1606_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6268_ (.A1(_1596_),
    .A2(_1602_),
    .B(_1606_),
    .ZN(_1607_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6269_ (.A1(\as2650.psl[1] ),
    .A2(_1195_),
    .ZN(_1608_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6270_ (.A1(_1607_),
    .A2(_1608_),
    .Z(_1609_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6271_ (.A1(_1590_),
    .A2(_1609_),
    .ZN(_1610_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _6272_ (.A1(_0608_),
    .A2(_0758_),
    .A3(_0854_),
    .A4(_1600_),
    .ZN(_1611_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6273_ (.A1(_1596_),
    .A2(_1611_),
    .ZN(_1612_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _6274_ (.A1(_1590_),
    .A2(_1209_),
    .A3(_1594_),
    .B1(_1610_),
    .B2(_1612_),
    .ZN(_1613_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6275_ (.I(_0320_),
    .Z(_1614_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6276_ (.A1(_1489_),
    .A2(_1614_),
    .ZN(_1615_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6277_ (.A1(_0876_),
    .A2(_0777_),
    .A3(_0662_),
    .ZN(_1616_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _6278_ (.A1(_1120_),
    .A2(_1087_),
    .A3(_1017_),
    .A4(_0949_),
    .ZN(_1617_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6279_ (.A1(_1616_),
    .A2(_1617_),
    .B(_1210_),
    .ZN(_1618_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6280_ (.I(_4081_),
    .Z(_1619_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6281_ (.A1(_1619_),
    .A2(_0373_),
    .ZN(_1620_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6282_ (.A1(_0373_),
    .A2(_1618_),
    .B1(_1620_),
    .B2(_1225_),
    .ZN(_1621_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6283_ (.I(_0552_),
    .Z(_1622_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6284_ (.A1(_4329_),
    .A2(_1459_),
    .ZN(_1623_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6285_ (.A1(_0487_),
    .A2(_1623_),
    .B(_1462_),
    .C(_4371_),
    .ZN(_1624_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _6286_ (.A1(_1622_),
    .A2(_1496_),
    .B(_1520_),
    .C(_1624_),
    .ZN(_1625_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6287_ (.I(_0546_),
    .Z(_1626_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _6288_ (.A1(_4320_),
    .A2(_4399_),
    .A3(_0564_),
    .B(_1478_),
    .ZN(_1627_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6289_ (.A1(_1524_),
    .A2(_1626_),
    .B(_1627_),
    .ZN(_1628_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _6290_ (.A1(_4449_),
    .A2(_1468_),
    .A3(_0481_),
    .ZN(_1629_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _6291_ (.A1(_0736_),
    .A2(_0738_),
    .B(_1629_),
    .ZN(_1630_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6292_ (.A1(_4049_),
    .A2(_0503_),
    .B(_1630_),
    .ZN(_1631_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6293_ (.A1(_1465_),
    .A2(_0476_),
    .ZN(_1632_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6294_ (.I(_1632_),
    .Z(_1633_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6295_ (.A1(_1633_),
    .A2(_1622_),
    .A3(_1469_),
    .ZN(_1634_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6296_ (.A1(_4319_),
    .A2(_1459_),
    .ZN(_1635_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6297_ (.A1(_1473_),
    .A2(_0483_),
    .ZN(_1636_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6298_ (.A1(_1634_),
    .A2(_1635_),
    .A3(_1636_),
    .ZN(_1637_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _6299_ (.A1(_4359_),
    .A2(_0448_),
    .A3(_0290_),
    .ZN(_1638_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6300_ (.I(_0677_),
    .Z(_1639_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6301_ (.A1(_4371_),
    .A2(_1639_),
    .ZN(_1640_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _6302_ (.A1(_0446_),
    .A2(_1495_),
    .A3(_1638_),
    .A4(_1640_),
    .ZN(_1641_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _6303_ (.A1(_0369_),
    .A2(_0363_),
    .A3(_0364_),
    .A4(_0372_),
    .ZN(_1642_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6304_ (.I(_1265_),
    .Z(_1643_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6305_ (.A1(_1643_),
    .A2(_0731_),
    .ZN(_1644_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6306_ (.A1(_1473_),
    .A2(_1644_),
    .B(_1515_),
    .ZN(_1645_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _6307_ (.A1(_0490_),
    .A2(_1641_),
    .B1(_1642_),
    .B2(_0302_),
    .C(_1645_),
    .ZN(_1646_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _6308_ (.A1(_1628_),
    .A2(_1631_),
    .A3(_1637_),
    .A4(_1646_),
    .ZN(_1647_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6309_ (.A1(_1625_),
    .A2(_1647_),
    .Z(_1648_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6310_ (.A1(_0666_),
    .A2(_0448_),
    .ZN(_1649_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6311_ (.I(_1649_),
    .Z(_1650_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6312_ (.A1(_1650_),
    .A2(_0673_),
    .ZN(_1651_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6313_ (.A1(_1122_),
    .A2(_0475_),
    .ZN(_1652_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6314_ (.A1(_0475_),
    .A2(_1618_),
    .B(_1652_),
    .C(_1524_),
    .ZN(_1653_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6315_ (.I(_1465_),
    .Z(_1654_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6316_ (.A1(_0813_),
    .A2(_1468_),
    .A3(_0496_),
    .ZN(_1655_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6317_ (.I(net2),
    .ZN(_1656_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6318_ (.I(_1656_),
    .Z(_1657_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6319_ (.I(_1657_),
    .Z(_1658_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6320_ (.I(_1658_),
    .Z(_1659_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6321_ (.I(\as2650.psl[6] ),
    .Z(_1660_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6322_ (.A1(_1660_),
    .A2(_1658_),
    .ZN(_1661_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6323_ (.A1(_0476_),
    .A2(_1659_),
    .B(_1661_),
    .ZN(_1662_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _6324_ (.A1(_1654_),
    .A2(_4370_),
    .A3(_1655_),
    .A4(_1662_),
    .ZN(_1663_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6325_ (.A1(_1650_),
    .A2(_1653_),
    .A3(_1663_),
    .ZN(_1664_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6326_ (.A1(_1090_),
    .A2(_1650_),
    .B(_0793_),
    .C(_1664_),
    .ZN(_1665_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6327_ (.A1(_4180_),
    .A2(_1651_),
    .B(_1665_),
    .ZN(_1666_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6328_ (.A1(_1561_),
    .A2(_1099_),
    .A3(_4199_),
    .ZN(_1667_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6329_ (.I(_4185_),
    .Z(_1668_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _6330_ (.A1(_1619_),
    .A2(_4156_),
    .A3(_1667_),
    .A4(_1668_),
    .ZN(_1669_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6331_ (.I(_4318_),
    .Z(_1670_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _6332_ (.A1(_0793_),
    .A2(_1213_),
    .A3(_1669_),
    .B(_1670_),
    .ZN(_1671_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6333_ (.I(_1023_),
    .Z(_1672_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6334_ (.I(_1143_),
    .Z(_1673_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6335_ (.I(_1673_),
    .Z(_1674_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6336_ (.A1(_1672_),
    .A2(_1095_),
    .A3(_1674_),
    .ZN(_1675_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6337_ (.I(_0676_),
    .Z(_1676_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6338_ (.I(_0787_),
    .Z(_1677_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6339_ (.I(_0883_),
    .Z(_1678_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6340_ (.I(_0953_),
    .Z(_1679_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6341_ (.I(_1679_),
    .Z(_1680_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _6342_ (.A1(_1676_),
    .A2(_1677_),
    .A3(_1678_),
    .A4(_1680_),
    .ZN(_1681_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6343_ (.A1(_1675_),
    .A2(_1681_),
    .B(_0412_),
    .ZN(_1682_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _6344_ (.A1(_1666_),
    .A2(_1671_),
    .B1(_1682_),
    .B2(_1670_),
    .C(_0386_),
    .ZN(_1683_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6345_ (.A1(_1615_),
    .A2(_1621_),
    .B(_1648_),
    .C(_1683_),
    .ZN(_1684_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6346_ (.A1(_1589_),
    .A2(_1613_),
    .B(_1684_),
    .ZN(_1685_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6347_ (.I(_0350_),
    .Z(_1686_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6348_ (.I(_1686_),
    .Z(_1687_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6349_ (.A1(_1660_),
    .A2(_1648_),
    .B(_1687_),
    .ZN(_1688_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6350_ (.A1(_1685_),
    .A2(_1688_),
    .ZN(_0093_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6351_ (.I(_1686_),
    .Z(_1689_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6352_ (.I(\as2650.psl[7] ),
    .Z(_1690_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6353_ (.I(_4402_),
    .Z(_1691_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6354_ (.I(_4414_),
    .Z(_1692_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6355_ (.I(_1692_),
    .Z(_1693_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6356_ (.I(_1693_),
    .Z(_1694_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6357_ (.I(_1639_),
    .Z(_1695_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6358_ (.A1(_4450_),
    .A2(_4306_),
    .ZN(_1696_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6359_ (.I(_1696_),
    .Z(_1697_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6360_ (.I(_0520_),
    .Z(_1698_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6361_ (.A1(_1668_),
    .A2(_1697_),
    .B1(_1698_),
    .B2(_1213_),
    .ZN(_1699_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6362_ (.I(_4306_),
    .Z(_1700_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6363_ (.I(_1700_),
    .Z(_1701_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _6364_ (.A1(_4414_),
    .A2(_0672_),
    .B1(_1561_),
    .B2(_1094_),
    .C1(_4189_),
    .C2(_1022_),
    .ZN(_1702_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _6365_ (.A1(_0882_),
    .A2(_4192_),
    .B1(_1089_),
    .B2(_1143_),
    .C1(_4215_),
    .C2(_0675_),
    .ZN(_1703_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6366_ (.A1(_4387_),
    .A2(_0620_),
    .ZN(_1704_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6367_ (.A1(_4372_),
    .A2(_1467_),
    .A3(_1704_),
    .ZN(_1705_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6368_ (.A1(_1679_),
    .A2(_4207_),
    .B1(_4209_),
    .B2(_0786_),
    .C(_1705_),
    .ZN(_1706_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _6369_ (.A1(_1702_),
    .A2(_1703_),
    .A3(_1706_),
    .Z(_1707_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _6370_ (.I(_0675_),
    .ZN(_1708_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6371_ (.I(net10),
    .ZN(_1709_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6372_ (.I(_1709_),
    .Z(_1710_));
 gf180mcu_fd_sc_mcu7t5v0__oai222_1 _6373_ (.A1(\as2650.psl[7] ),
    .A2(_1214_),
    .B1(_1708_),
    .B2(_0610_),
    .C1(_0609_),
    .C2(_1710_),
    .ZN(_1711_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _6374_ (.I(_0784_),
    .ZN(_1712_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6375_ (.I(_1712_),
    .Z(_1713_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6376_ (.A1(_0549_),
    .A2(_1021_),
    .ZN(_1714_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _6377_ (.A1(\as2650.psl[1] ),
    .A2(_1713_),
    .B1(_1658_),
    .B2(_1660_),
    .C(_1714_),
    .ZN(_1715_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6378_ (.I(_0881_),
    .ZN(_1716_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6379_ (.I(_1716_),
    .Z(_1717_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6380_ (.I(_1717_),
    .Z(_1718_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6381_ (.A1(\as2650.overflow ),
    .A2(_1718_),
    .B1(_1500_),
    .B2(\as2650.psl[5] ),
    .ZN(_1719_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _6382_ (.A1(_1711_),
    .A2(_1715_),
    .A3(_1719_),
    .Z(_1720_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6383_ (.A1(_1654_),
    .A2(_1720_),
    .B(_1704_),
    .C(_1467_),
    .ZN(_1721_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6384_ (.A1(_1465_),
    .A2(_1467_),
    .ZN(_1722_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6385_ (.I(\as2650.psu[4] ),
    .ZN(_1723_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6386_ (.A1(_0699_),
    .A2(_1708_),
    .B1(_1709_),
    .B2(\as2650.psu[3] ),
    .ZN(_1724_));
 gf180mcu_fd_sc_mcu7t5v0__oai222_1 _6387_ (.A1(_0708_),
    .A2(_1712_),
    .B1(_1718_),
    .B2(\as2650.psu[2] ),
    .C1(\as2650.psu[7] ),
    .C2(_1214_),
    .ZN(_1725_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6388_ (.A1(_1723_),
    .A2(_1021_),
    .B(_1724_),
    .C(_1725_),
    .ZN(_1726_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _6389_ (.A1(\as2650.psu[5] ),
    .A2(_1501_),
    .B1(_1658_),
    .B2(net28),
    .C(_1726_),
    .ZN(_1727_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _6390_ (.A1(_4388_),
    .A2(_0621_),
    .A3(_1722_),
    .A4(_1727_),
    .ZN(_1728_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6391_ (.I(_4248_),
    .Z(_1729_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6392_ (.A1(_1729_),
    .A2(_1469_),
    .ZN(_1730_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6393_ (.A1(_1707_),
    .A2(_1721_),
    .B(_1728_),
    .C(_1730_),
    .ZN(_1731_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6394_ (.A1(_0477_),
    .A2(_1494_),
    .ZN(_1732_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6395_ (.A1(_1690_),
    .A2(_0410_),
    .A3(_1730_),
    .ZN(_1733_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6396_ (.A1(_1732_),
    .A2(_1733_),
    .ZN(_1734_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6397_ (.A1(_1692_),
    .A2(_1476_),
    .ZN(_1735_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6398_ (.A1(_1731_),
    .A2(_1734_),
    .B1(_1735_),
    .B2(_1690_),
    .ZN(_1736_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6399_ (.A1(_1210_),
    .A2(_1524_),
    .ZN(_1737_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6400_ (.A1(_1479_),
    .A2(_1736_),
    .B(_1737_),
    .ZN(_1738_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6401_ (.A1(_1701_),
    .A2(_1738_),
    .ZN(_1739_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6402_ (.A1(_1699_),
    .A2(_1739_),
    .B(_1639_),
    .ZN(_1740_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6403_ (.A1(_1694_),
    .A2(_1695_),
    .B(_1740_),
    .ZN(_1741_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6404_ (.A1(_1590_),
    .A2(_1208_),
    .B(_1610_),
    .C(_4050_),
    .ZN(_1742_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6405_ (.A1(_1474_),
    .A2(_0371_),
    .ZN(_1743_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6406_ (.A1(_1614_),
    .A2(_1737_),
    .A3(_1743_),
    .ZN(_1744_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6407_ (.A1(_1619_),
    .A2(_0373_),
    .B(_1744_),
    .ZN(_1745_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6408_ (.A1(_1691_),
    .A2(_1741_),
    .B1(_1742_),
    .B2(_1745_),
    .ZN(_1746_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6409_ (.I0(_1690_),
    .I1(_1746_),
    .S(_1648_),
    .Z(_1747_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6410_ (.A1(_1689_),
    .A2(_1747_),
    .Z(_1748_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6411_ (.I(_1748_),
    .Z(_0094_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6412_ (.A1(_0337_),
    .A2(_0348_),
    .ZN(_1749_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6413_ (.A1(_4364_),
    .A2(_1749_),
    .Z(_1750_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6414_ (.I(_1750_),
    .Z(_1751_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6415_ (.I(_1676_),
    .Z(_1752_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6416_ (.A1(_0342_),
    .A2(_1752_),
    .ZN(_1753_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6417_ (.I(_1750_),
    .Z(_1754_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6418_ (.A1(_0736_),
    .A2(_1215_),
    .ZN(_1755_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6419_ (.A1(_0397_),
    .A2(_1755_),
    .ZN(_1756_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _6420_ (.A1(_0339_),
    .A2(_4246_),
    .A3(_4256_),
    .A4(_1756_),
    .ZN(_1757_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6421_ (.A1(_1754_),
    .A2(_1757_),
    .ZN(_1758_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6422_ (.I(_1758_),
    .Z(_1759_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6423_ (.A1(_1751_),
    .A2(_1753_),
    .B1(_1759_),
    .B2(_4372_),
    .ZN(_0095_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6424_ (.A1(_0342_),
    .A2(_1677_),
    .ZN(_1760_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6425_ (.I(_1754_),
    .Z(_1761_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6426_ (.A1(_0476_),
    .A2(_1759_),
    .B1(_1760_),
    .B2(_1761_),
    .ZN(_0096_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6427_ (.A1(_1678_),
    .A2(_1751_),
    .B1(_1759_),
    .B2(_0437_),
    .ZN(_1762_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6428_ (.I(_1762_),
    .ZN(_0097_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6429_ (.A1(_4341_),
    .A2(_1245_),
    .ZN(_1763_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6430_ (.I(_1763_),
    .Z(_1764_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6431_ (.A1(_0348_),
    .A2(_1502_),
    .ZN(_1765_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6432_ (.A1(_0348_),
    .A2(_1764_),
    .B(_1765_),
    .ZN(_1766_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6433_ (.A1(_0615_),
    .A2(_1761_),
    .B1(_1759_),
    .B2(_1766_),
    .ZN(_0098_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6434_ (.A1(_1674_),
    .A2(_1751_),
    .B1(_1758_),
    .B2(_0494_),
    .ZN(_1767_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6435_ (.I(_1767_),
    .ZN(_0099_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6436_ (.A1(_0413_),
    .A2(_1751_),
    .B1(_1758_),
    .B2(_0666_),
    .ZN(_1768_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6437_ (.I(_1768_),
    .ZN(_0100_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _6438_ (.A1(_0700_),
    .A2(_1348_),
    .A3(_1351_),
    .A4(_1367_),
    .ZN(_1769_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6439_ (.I(_1769_),
    .Z(_1770_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6440_ (.I(_1770_),
    .Z(_1771_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6441_ (.I(_1770_),
    .Z(_1772_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6442_ (.A1(\as2650.stack[0][8] ),
    .A2(_1772_),
    .ZN(_1773_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6443_ (.A1(_1386_),
    .A2(_1771_),
    .B(_1773_),
    .ZN(_0101_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6444_ (.I(_1769_),
    .Z(_1774_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6445_ (.A1(\as2650.stack[0][9] ),
    .A2(_1774_),
    .ZN(_1775_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6446_ (.A1(_1396_),
    .A2(_1771_),
    .B(_1775_),
    .ZN(_0102_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6447_ (.A1(\as2650.stack[0][10] ),
    .A2(_1774_),
    .ZN(_1776_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6448_ (.A1(_1404_),
    .A2(_1771_),
    .B(_1776_),
    .ZN(_0103_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6449_ (.A1(\as2650.stack[0][11] ),
    .A2(_1774_),
    .ZN(_1777_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6450_ (.A1(_1414_),
    .A2(_1771_),
    .B(_1777_),
    .ZN(_0104_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6451_ (.A1(\as2650.stack[0][12] ),
    .A2(_1774_),
    .ZN(_1778_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6452_ (.A1(_1420_),
    .A2(_1772_),
    .B(_1778_),
    .ZN(_0105_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6453_ (.A1(\as2650.stack[0][13] ),
    .A2(_1770_),
    .ZN(_1779_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6454_ (.A1(_1427_),
    .A2(_1772_),
    .B(_1779_),
    .ZN(_0106_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6455_ (.A1(\as2650.stack[0][14] ),
    .A2(_1770_),
    .ZN(_1780_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6456_ (.A1(_1434_),
    .A2(_1772_),
    .B(_1780_),
    .ZN(_0107_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6457_ (.I(_1385_),
    .Z(_1781_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6458_ (.I(_1268_),
    .Z(_1782_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6459_ (.A1(_1348_),
    .A2(_1366_),
    .ZN(_1783_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6460_ (.A1(_1346_),
    .A2(_1782_),
    .A3(_1783_),
    .ZN(_1784_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6461_ (.I(_1784_),
    .Z(_1785_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6462_ (.I(_1785_),
    .Z(_1786_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6463_ (.I(_1785_),
    .Z(_1787_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6464_ (.A1(\as2650.stack[6][8] ),
    .A2(_1787_),
    .ZN(_1788_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6465_ (.A1(_1781_),
    .A2(_1786_),
    .B(_1788_),
    .ZN(_0108_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6466_ (.I(_1395_),
    .Z(_1789_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6467_ (.I(_1784_),
    .Z(_1790_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6468_ (.A1(\as2650.stack[6][9] ),
    .A2(_1790_),
    .ZN(_1791_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6469_ (.A1(_1789_),
    .A2(_1786_),
    .B(_1791_),
    .ZN(_0109_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6470_ (.I(_1403_),
    .Z(_1792_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6471_ (.A1(\as2650.stack[6][10] ),
    .A2(_1790_),
    .ZN(_1793_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6472_ (.A1(_1792_),
    .A2(_1786_),
    .B(_1793_),
    .ZN(_0110_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6473_ (.I(_1413_),
    .Z(_1794_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6474_ (.A1(\as2650.stack[6][11] ),
    .A2(_1790_),
    .ZN(_1795_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6475_ (.A1(_1794_),
    .A2(_1786_),
    .B(_1795_),
    .ZN(_0111_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6476_ (.I(_1419_),
    .Z(_1796_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6477_ (.A1(\as2650.stack[6][12] ),
    .A2(_1790_),
    .ZN(_1797_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6478_ (.A1(_1796_),
    .A2(_1787_),
    .B(_1797_),
    .ZN(_0112_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6479_ (.I(_1426_),
    .Z(_1798_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6480_ (.A1(\as2650.stack[6][13] ),
    .A2(_1785_),
    .ZN(_1799_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6481_ (.A1(_1798_),
    .A2(_1787_),
    .B(_1799_),
    .ZN(_0113_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6482_ (.I(_1433_),
    .Z(_1800_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6483_ (.A1(\as2650.stack[6][14] ),
    .A2(_1785_),
    .ZN(_1801_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6484_ (.A1(_1800_),
    .A2(_1787_),
    .B(_1801_),
    .ZN(_0114_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6485_ (.A1(_0337_),
    .A2(_4245_),
    .ZN(_1802_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6486_ (.A1(_0524_),
    .A2(_4374_),
    .ZN(_1803_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6487_ (.I(_1803_),
    .ZN(_1804_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _6488_ (.A1(_4413_),
    .A2(_1802_),
    .A3(_0536_),
    .A4(_1804_),
    .ZN(_1805_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6489_ (.I(_1805_),
    .Z(_1806_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6490_ (.A1(_4082_),
    .A2(_0516_),
    .ZN(_1807_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6491_ (.I(_1807_),
    .Z(_1808_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6492_ (.A1(_4357_),
    .A2(_4374_),
    .A3(_1808_),
    .ZN(_1809_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6493_ (.A1(_4293_),
    .A2(_0792_),
    .A3(_1809_),
    .ZN(_1810_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6494_ (.I(_1810_),
    .Z(_1811_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _6495_ (.A1(_0524_),
    .A2(_4310_),
    .A3(_0515_),
    .ZN(_1812_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6496_ (.A1(_0553_),
    .A2(_1812_),
    .ZN(_1813_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6497_ (.I(_1813_),
    .Z(_1814_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6498_ (.A1(_4356_),
    .A2(_1807_),
    .ZN(_1815_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6499_ (.A1(_4393_),
    .A2(_1815_),
    .ZN(_1816_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _6500_ (.A1(_0630_),
    .A2(_4307_),
    .A3(_1816_),
    .ZN(_1817_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6501_ (.I(_1817_),
    .Z(_1818_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6502_ (.A1(_0566_),
    .A2(_1808_),
    .ZN(_1819_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6503_ (.A1(_0367_),
    .A2(_0301_),
    .A3(_1816_),
    .ZN(_1820_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6504_ (.I(_1820_),
    .Z(_1821_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6505_ (.A1(_1818_),
    .A2(_1819_),
    .A3(_1821_),
    .ZN(_1822_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6506_ (.A1(\as2650.cycle[9] ),
    .A2(_4281_),
    .ZN(_1823_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _6507_ (.A1(_4284_),
    .A2(_0419_),
    .A3(_1803_),
    .A4(_1823_),
    .ZN(_1824_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6508_ (.A1(_0543_),
    .A2(_1260_),
    .A3(_1824_),
    .ZN(_1825_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _6509_ (.I(_1825_),
    .ZN(_1826_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _6510_ (.A1(_1811_),
    .A2(_1814_),
    .A3(_1822_),
    .A4(_1826_),
    .ZN(_1827_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _6511_ (.A1(_0549_),
    .A2(_0559_),
    .B(_1806_),
    .C(_1827_),
    .ZN(_1828_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6512_ (.I(_1828_),
    .Z(_1829_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6513_ (.A1(_1729_),
    .A2(_1829_),
    .ZN(_1830_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6514_ (.I(_1830_),
    .Z(_1831_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6515_ (.I(_1831_),
    .Z(_1832_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6516_ (.I(_1825_),
    .Z(_1833_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6517_ (.I(_1833_),
    .Z(_1834_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6518_ (.I(_1805_),
    .Z(_1835_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6519_ (.I(_1820_),
    .Z(_1836_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6520_ (.I(_1813_),
    .Z(_1837_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6521_ (.A1(_0676_),
    .A2(_1837_),
    .ZN(_1838_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6522_ (.A1(_4158_),
    .A2(_4215_),
    .Z(_1839_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6523_ (.A1(_0680_),
    .A2(_1808_),
    .ZN(_1840_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6524_ (.A1(_1839_),
    .A2(_1840_),
    .B(_1810_),
    .ZN(_1841_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _6525_ (.A1(_4449_),
    .A2(_0546_),
    .A3(_1809_),
    .ZN(_1842_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6526_ (.A1(_0674_),
    .A2(_1811_),
    .B1(_1838_),
    .B2(_1841_),
    .C(_1842_),
    .ZN(_1843_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6527_ (.A1(_0673_),
    .A2(_1842_),
    .ZN(_1844_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6528_ (.A1(_1821_),
    .A2(_1844_),
    .ZN(_1845_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6529_ (.A1(_0662_),
    .A2(_1836_),
    .B1(_1843_),
    .B2(_1845_),
    .ZN(_1846_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6530_ (.A1(_1806_),
    .A2(_1846_),
    .ZN(_1847_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6531_ (.A1(_0659_),
    .A2(_1835_),
    .B(_1833_),
    .C(_1847_),
    .ZN(_1848_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6532_ (.A1(_0651_),
    .A2(_1834_),
    .B(_1848_),
    .ZN(_1849_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6533_ (.I(_1819_),
    .Z(_1850_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6534_ (.I0(_0638_),
    .I1(_1849_),
    .S(_1850_),
    .Z(_1851_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6535_ (.I(_1851_),
    .ZN(_1852_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6536_ (.A1(_0740_),
    .A2(_1812_),
    .ZN(_1853_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6537_ (.I(_1853_),
    .Z(_1854_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6538_ (.A1(_1729_),
    .A2(_1829_),
    .B(_1854_),
    .C(_0322_),
    .ZN(_1855_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6539_ (.I(_1855_),
    .Z(_1856_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6540_ (.I0(\as2650.r123[0][5] ),
    .I1(\as2650.r123_2[0][5] ),
    .S(\as2650.psl[4] ),
    .Z(_1857_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6541_ (.I(_1857_),
    .Z(_1858_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6542_ (.I(_1858_),
    .Z(_1859_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6543_ (.I0(\as2650.r123[0][4] ),
    .I1(\as2650.r123_2[0][4] ),
    .S(_4088_),
    .Z(_1860_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6544_ (.I(_1860_),
    .Z(_1861_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _6545_ (.A1(_4149_),
    .A2(_4159_),
    .A3(_1859_),
    .A4(_1861_),
    .Z(_1862_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6546_ (.I(_1862_),
    .Z(_1863_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6547_ (.I(_1859_),
    .Z(_1864_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6548_ (.I(_1861_),
    .Z(_1865_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6549_ (.A1(_4160_),
    .A2(_1864_),
    .B1(_1865_),
    .B2(_0752_),
    .ZN(_1866_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6550_ (.A1(_1863_),
    .A2(_1866_),
    .ZN(_1867_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6551_ (.I0(\as2650.r123[0][0] ),
    .I1(\as2650.r123_2[0][0] ),
    .S(_4061_),
    .Z(_1868_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6552_ (.I(_1868_),
    .Z(_1869_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6553_ (.A1(_4105_),
    .A2(_1869_),
    .ZN(_1870_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6554_ (.I0(\as2650.r123[0][1] ),
    .I1(\as2650.r123_2[0][1] ),
    .S(_4088_),
    .Z(_1871_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6555_ (.I(_1871_),
    .Z(_1872_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6556_ (.A1(_4117_),
    .A2(_1872_),
    .ZN(_1873_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6557_ (.I0(\as2650.r123[0][3] ),
    .I1(\as2650.r123_2[0][3] ),
    .S(_4088_),
    .Z(_1874_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6558_ (.I(_1874_),
    .Z(_1875_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6559_ (.A1(_4138_),
    .A2(_1875_),
    .ZN(_1876_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _6560_ (.A1(_1870_),
    .A2(_1873_),
    .A3(_1876_),
    .Z(_1877_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6561_ (.A1(_1867_),
    .A2(_1877_),
    .ZN(_1878_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6562_ (.A1(_0589_),
    .A2(_1865_),
    .ZN(_1879_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6563_ (.A1(_4118_),
    .A2(_1869_),
    .Z(_1880_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6564_ (.A1(_4127_),
    .A2(_1872_),
    .ZN(_1881_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6565_ (.I(_1875_),
    .Z(_1882_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6566_ (.A1(_4150_),
    .A2(_1882_),
    .ZN(_1883_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _6567_ (.A1(_1880_),
    .A2(_1881_),
    .A3(_1883_),
    .ZN(_1884_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6568_ (.A1(_1879_),
    .A2(_1884_),
    .ZN(_1885_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6569_ (.A1(_1881_),
    .A2(_1883_),
    .ZN(_1886_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6570_ (.A1(_1881_),
    .A2(_1883_),
    .ZN(_1887_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6571_ (.A1(_1880_),
    .A2(_1886_),
    .B(_1887_),
    .ZN(_1888_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6572_ (.I0(\as2650.r123[0][2] ),
    .I1(\as2650.r123_2[0][2] ),
    .S(_4108_),
    .Z(_1889_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6573_ (.I(_1889_),
    .Z(_1890_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6574_ (.A1(_0918_),
    .A2(_1890_),
    .ZN(_1891_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6575_ (.A1(_1888_),
    .A2(_1891_),
    .ZN(_1892_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _6576_ (.A1(_1878_),
    .A2(_1885_),
    .A3(_1892_),
    .ZN(_1893_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6577_ (.A1(_1879_),
    .A2(_1884_),
    .ZN(_1894_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6578_ (.I(_1871_),
    .Z(_1895_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6579_ (.I(_1895_),
    .Z(_1896_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6580_ (.A1(_0588_),
    .A2(_1896_),
    .ZN(_1897_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6581_ (.I(_1869_),
    .Z(_1898_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6582_ (.A1(_4128_),
    .A2(_1898_),
    .ZN(_1899_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6583_ (.A1(_0588_),
    .A2(_1882_),
    .B1(_1896_),
    .B2(_4139_),
    .ZN(_1900_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6584_ (.A1(_1876_),
    .A2(_1897_),
    .B1(_1899_),
    .B2(_1900_),
    .ZN(_1901_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6585_ (.I(_1890_),
    .Z(_1902_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6586_ (.A1(_0844_),
    .A2(_1902_),
    .ZN(_1903_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6587_ (.A1(_1901_),
    .A2(_1903_),
    .Z(_1904_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6588_ (.I(_1902_),
    .Z(_1905_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6589_ (.I(_1905_),
    .Z(_1906_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6590_ (.A1(_0876_),
    .A2(_1906_),
    .A3(_1901_),
    .ZN(_1907_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6591_ (.A1(_1894_),
    .A2(_1904_),
    .B(_1907_),
    .ZN(_1908_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6592_ (.A1(_1893_),
    .A2(_1908_),
    .Z(_1909_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _6593_ (.A1(_0844_),
    .A2(_0752_),
    .A3(_1896_),
    .A4(_1898_),
    .Z(_1910_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6594_ (.A1(_0776_),
    .A2(_1902_),
    .Z(_1911_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6595_ (.A1(_1905_),
    .A2(_1910_),
    .ZN(_1912_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6596_ (.A1(_1910_),
    .A2(_1911_),
    .B(_1912_),
    .ZN(_1913_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6597_ (.A1(_4139_),
    .A2(_1895_),
    .ZN(_1914_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6598_ (.I(_1882_),
    .Z(_1915_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6599_ (.A1(_0588_),
    .A2(_1915_),
    .ZN(_1916_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _6600_ (.A1(_1914_),
    .A2(_1916_),
    .A3(_1899_),
    .Z(_1917_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6601_ (.A1(_1913_),
    .A2(_1917_),
    .B(_1912_),
    .ZN(_1918_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6602_ (.A1(_1894_),
    .A2(_1904_),
    .Z(_1919_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6603_ (.A1(_1918_),
    .A2(_1919_),
    .ZN(_1920_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6604_ (.A1(_1918_),
    .A2(_1919_),
    .Z(_1921_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6605_ (.I(_1896_),
    .Z(_1922_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6606_ (.I(_1898_),
    .Z(_1923_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6607_ (.A1(_0601_),
    .A2(_1923_),
    .Z(_1924_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _6608_ (.A1(_0777_),
    .A2(_1906_),
    .A3(_1922_),
    .A4(_1924_),
    .Z(_1925_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6609_ (.A1(_0601_),
    .A2(_1905_),
    .ZN(_1926_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _6610_ (.A1(_0776_),
    .A2(_0589_),
    .A3(_1922_),
    .A4(_1898_),
    .ZN(_1927_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6611_ (.I0(_1905_),
    .I1(_1926_),
    .S(_1927_),
    .Z(_1928_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6612_ (.A1(_0776_),
    .A2(_1922_),
    .B1(_1923_),
    .B2(_0876_),
    .ZN(_1929_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6613_ (.A1(_1910_),
    .A2(_1929_),
    .Z(_1930_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6614_ (.A1(_1928_),
    .A2(_1930_),
    .ZN(_1931_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6615_ (.A1(_1925_),
    .A2(_1931_),
    .ZN(_1932_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6616_ (.A1(_1913_),
    .A2(_1917_),
    .ZN(_1933_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6617_ (.A1(_1932_),
    .A2(_1933_),
    .ZN(_1934_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6618_ (.A1(_1921_),
    .A2(_1934_),
    .ZN(_1935_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6619_ (.A1(_1893_),
    .A2(_1908_),
    .ZN(_1936_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6620_ (.A1(_1920_),
    .A2(_1935_),
    .B(_1936_),
    .ZN(_1937_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6621_ (.A1(_1888_),
    .A2(_1891_),
    .Z(_1938_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6622_ (.A1(_1878_),
    .A2(_1885_),
    .ZN(_1939_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6623_ (.A1(_1878_),
    .A2(_1885_),
    .ZN(_1940_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6624_ (.A1(_1939_),
    .A2(_1892_),
    .B(_1940_),
    .ZN(_1941_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6625_ (.A1(_4117_),
    .A2(_1874_),
    .ZN(_1942_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6626_ (.A1(_1873_),
    .A2(_1876_),
    .Z(_1943_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6627_ (.A1(_1942_),
    .A2(_1914_),
    .B1(_1943_),
    .B2(_1870_),
    .ZN(_1944_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6628_ (.A1(_4118_),
    .A2(_1890_),
    .ZN(_1945_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6629_ (.A1(_1944_),
    .A2(_1945_),
    .Z(_1946_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _6630_ (.A1(_1863_),
    .A2(_1866_),
    .A3(_1877_),
    .Z(_1947_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6631_ (.A1(\as2650.r0[1] ),
    .A2(_1857_),
    .ZN(_1948_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6632_ (.A1(\as2650.r0[2] ),
    .A2(_1860_),
    .ZN(_1949_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6633_ (.A1(\as2650.r0[0] ),
    .A2(_4090_),
    .ZN(_1950_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _6634_ (.A1(_1948_),
    .A2(_1949_),
    .A3(_1950_),
    .ZN(_1951_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6635_ (.A1(_4127_),
    .A2(_1874_),
    .ZN(_1952_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6636_ (.A1(\as2650.r0[6] ),
    .A2(_1868_),
    .ZN(_1953_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6637_ (.A1(_4105_),
    .A2(_1895_),
    .ZN(_1954_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _6638_ (.A1(_1952_),
    .A2(_1953_),
    .A3(_1954_),
    .ZN(_1955_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _6639_ (.A1(_1862_),
    .A2(_1951_),
    .A3(_1955_),
    .ZN(_1956_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6640_ (.A1(_1947_),
    .A2(_1956_),
    .ZN(_1957_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6641_ (.A1(_1946_),
    .A2(_1957_),
    .Z(_1958_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6642_ (.A1(_1941_),
    .A2(_1958_),
    .ZN(_1959_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6643_ (.A1(_1938_),
    .A2(_1959_),
    .Z(_1960_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6644_ (.A1(_1909_),
    .A2(_1937_),
    .B(_1960_),
    .ZN(_1961_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6645_ (.A1(_1941_),
    .A2(_1958_),
    .ZN(_1962_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6646_ (.A1(_1938_),
    .A2(_1959_),
    .B(_1962_),
    .ZN(_1963_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6647_ (.A1(_0988_),
    .A2(_1906_),
    .A3(_1944_),
    .ZN(_1964_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6648_ (.A1(_1947_),
    .A2(_1956_),
    .Z(_1965_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6649_ (.A1(_1946_),
    .A2(_1957_),
    .B(_1965_),
    .ZN(_1966_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6650_ (.A1(_4105_),
    .A2(_1889_),
    .ZN(_1967_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6651_ (.I(\as2650.r0[5] ),
    .Z(_1968_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6652_ (.A1(_1968_),
    .A2(_1875_),
    .ZN(_1969_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6653_ (.A1(_4128_),
    .A2(_1874_),
    .B1(_1872_),
    .B2(_1968_),
    .ZN(_1970_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6654_ (.A1(_1881_),
    .A2(_1969_),
    .B1(_1970_),
    .B2(_1953_),
    .ZN(_1971_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6655_ (.A1(_4061_),
    .A2(\as2650.r123_2[0][7] ),
    .ZN(_1972_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6656_ (.A1(_4108_),
    .A2(_1182_),
    .B(_1972_),
    .ZN(_1973_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6657_ (.A1(_4159_),
    .A2(_1973_),
    .ZN(_1974_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6658_ (.A1(_1971_),
    .A2(_1974_),
    .ZN(_1975_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6659_ (.A1(_1967_),
    .A2(_1975_),
    .Z(_1976_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6660_ (.A1(_1863_),
    .A2(_1951_),
    .ZN(_1977_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6661_ (.I(_1955_),
    .ZN(_1978_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6662_ (.A1(_1863_),
    .A2(_1951_),
    .ZN(_1979_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6663_ (.A1(_1977_),
    .A2(_1978_),
    .B(_1979_),
    .ZN(_1980_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6664_ (.A1(_4098_),
    .A2(_1872_),
    .ZN(_1981_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6665_ (.A1(\as2650.r0[7] ),
    .A2(_1869_),
    .ZN(_1982_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _6666_ (.A1(_1942_),
    .A2(_1981_),
    .A3(_1982_),
    .Z(_1983_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6667_ (.A1(_4160_),
    .A2(_1859_),
    .ZN(_1984_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6668_ (.A1(\as2650.r0[1] ),
    .A2(_4089_),
    .ZN(_1985_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6669_ (.A1(_4149_),
    .A2(_1858_),
    .B1(_4091_),
    .B2(_4159_),
    .ZN(_1986_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6670_ (.A1(_1984_),
    .A2(_1985_),
    .B1(_1986_),
    .B2(_1949_),
    .ZN(_1987_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6671_ (.A1(\as2650.r0[3] ),
    .A2(_1860_),
    .ZN(_1988_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6672_ (.A1(\as2650.r0[2] ),
    .A2(_1858_),
    .ZN(_1989_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _6673_ (.A1(_1985_),
    .A2(_1988_),
    .A3(_1989_),
    .ZN(_1990_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6674_ (.A1(_1987_),
    .A2(_1990_),
    .ZN(_1991_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6675_ (.A1(_1983_),
    .A2(_1991_),
    .Z(_1992_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _6676_ (.A1(_1976_),
    .A2(_1980_),
    .A3(_1992_),
    .Z(_1993_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6677_ (.A1(_1966_),
    .A2(_1993_),
    .Z(_1994_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6678_ (.A1(_1964_),
    .A2(_1994_),
    .Z(_1995_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6679_ (.A1(_1963_),
    .A2(_1995_),
    .ZN(_1996_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6680_ (.A1(_1963_),
    .A2(_1995_),
    .ZN(_1997_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6681_ (.A1(_1961_),
    .A2(_1996_),
    .B(_1997_),
    .ZN(_1998_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6682_ (.I(_1966_),
    .ZN(_1999_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6683_ (.A1(_1999_),
    .A2(_1993_),
    .ZN(_2000_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6684_ (.A1(_1964_),
    .A2(_1994_),
    .ZN(_2001_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6685_ (.A1(_2000_),
    .A2(_2001_),
    .ZN(_2002_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6686_ (.I(_1973_),
    .Z(_2003_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6687_ (.A1(_0662_),
    .A2(_2003_),
    .A3(_1971_),
    .ZN(_2004_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6688_ (.I(_1906_),
    .Z(_2005_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6689_ (.A1(_4106_),
    .A2(_2005_),
    .A3(_1975_),
    .ZN(_2006_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6690_ (.A1(_2004_),
    .A2(_2006_),
    .ZN(_2007_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6691_ (.A1(_1980_),
    .A2(_1992_),
    .ZN(_2008_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6692_ (.A1(_1980_),
    .A2(_1992_),
    .ZN(_2009_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6693_ (.A1(_1976_),
    .A2(_2008_),
    .B(_2009_),
    .ZN(_2010_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6694_ (.A1(_4099_),
    .A2(_1890_),
    .ZN(_2011_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6695_ (.A1(_4098_),
    .A2(_1875_),
    .ZN(_2012_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6696_ (.A1(_1942_),
    .A2(_1981_),
    .Z(_2013_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6697_ (.A1(_1873_),
    .A2(_2012_),
    .B1(_2013_),
    .B2(_1982_),
    .ZN(_2014_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6698_ (.A1(_4150_),
    .A2(_1973_),
    .ZN(_2015_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6699_ (.A1(_2014_),
    .A2(_2015_),
    .ZN(_2016_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6700_ (.A1(_2011_),
    .A2(_2016_),
    .Z(_2017_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6701_ (.A1(_1987_),
    .A2(_1990_),
    .ZN(_2018_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6702_ (.A1(_1983_),
    .A2(_1991_),
    .B(_2018_),
    .ZN(_2019_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6703_ (.A1(_4075_),
    .A2(_1895_),
    .ZN(_2020_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6704_ (.A1(_4075_),
    .A2(_1882_),
    .ZN(_2021_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6705_ (.A1(_1954_),
    .A2(_2021_),
    .ZN(_2022_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6706_ (.A1(_1969_),
    .A2(_2020_),
    .B(_2022_),
    .ZN(_2023_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6707_ (.A1(\as2650.r0[2] ),
    .A2(_4090_),
    .ZN(_2024_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6708_ (.A1(_4138_),
    .A2(_1859_),
    .B1(_4091_),
    .B2(_4149_),
    .ZN(_2025_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6709_ (.A1(_1948_),
    .A2(_2024_),
    .B1(_2025_),
    .B2(_1988_),
    .ZN(_2026_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6710_ (.A1(_4127_),
    .A2(_1857_),
    .ZN(_2027_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6711_ (.A1(_4117_),
    .A2(_1861_),
    .Z(_2028_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _6712_ (.A1(_2024_),
    .A2(_2027_),
    .A3(_2028_),
    .Z(_2029_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6713_ (.A1(_2026_),
    .A2(_2029_),
    .Z(_2030_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6714_ (.A1(_2023_),
    .A2(_2030_),
    .Z(_2031_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _6715_ (.A1(_2017_),
    .A2(_2019_),
    .A3(_2031_),
    .ZN(_2032_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6716_ (.A1(_2010_),
    .A2(_2032_),
    .Z(_2033_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6717_ (.A1(_2007_),
    .A2(_2033_),
    .ZN(_2034_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6718_ (.A1(_2002_),
    .A2(_2034_),
    .Z(_2035_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6719_ (.A1(_1998_),
    .A2(_2035_),
    .Z(_2036_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6720_ (.I(_1853_),
    .Z(_2037_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6721_ (.I(_2037_),
    .Z(_2038_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6722_ (.A1(\as2650.r123_2[2][0] ),
    .A2(_1856_),
    .B1(_2036_),
    .B2(_2038_),
    .ZN(_2039_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6723_ (.A1(_1832_),
    .A2(_1852_),
    .B(_2039_),
    .ZN(_0115_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6724_ (.I(_1833_),
    .Z(_2040_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6725_ (.I(_1835_),
    .Z(_2041_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6726_ (.I(_1836_),
    .Z(_2042_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6727_ (.I(_1806_),
    .Z(_2043_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6728_ (.I(_1821_),
    .Z(_2044_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6729_ (.I(_1817_),
    .Z(_2045_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6730_ (.A1(_4253_),
    .A2(_0520_),
    .A3(_1816_),
    .ZN(_2046_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6731_ (.I(_2046_),
    .Z(_2047_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6732_ (.I(_2047_),
    .Z(_2048_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6733_ (.I(_1813_),
    .Z(_2049_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6734_ (.A1(_0786_),
    .A2(_2049_),
    .ZN(_2050_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6735_ (.A1(_4218_),
    .A2(_1837_),
    .B(_2050_),
    .C(_2047_),
    .ZN(_2051_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6736_ (.A1(_0791_),
    .A2(_2048_),
    .B(_1818_),
    .C(_2051_),
    .ZN(_2052_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6737_ (.A1(_0782_),
    .A2(_2045_),
    .B(_2052_),
    .ZN(_2053_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6738_ (.A1(_2044_),
    .A2(_2053_),
    .ZN(_2054_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6739_ (.A1(_0753_),
    .A2(_2042_),
    .B(_2043_),
    .C(_2054_),
    .ZN(_2055_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6740_ (.A1(_0802_),
    .A2(_2041_),
    .B(_1834_),
    .C(_2055_),
    .ZN(_2056_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6741_ (.I(_1850_),
    .Z(_2057_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6742_ (.A1(_0807_),
    .A2(_2040_),
    .B(_2056_),
    .C(_2057_),
    .ZN(_2058_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6743_ (.A1(_0565_),
    .A2(_1812_),
    .ZN(_2059_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6744_ (.A1(_0775_),
    .A2(_2059_),
    .ZN(_2060_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6745_ (.A1(_2058_),
    .A2(_2060_),
    .ZN(_2061_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6746_ (.A1(_2002_),
    .A2(_2034_),
    .ZN(_2062_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _6747_ (.A1(_1998_),
    .A2(_2035_),
    .B(_2062_),
    .ZN(_2063_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6748_ (.A1(_2010_),
    .A2(_2032_),
    .Z(_2064_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6749_ (.A1(_2007_),
    .A2(_2033_),
    .B(_2064_),
    .ZN(_2065_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6750_ (.A1(_0777_),
    .A2(_2003_),
    .A3(_2014_),
    .ZN(_2066_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6751_ (.A1(_1120_),
    .A2(_2005_),
    .A3(_2016_),
    .ZN(_2067_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6752_ (.A1(_2066_),
    .A2(_2067_),
    .ZN(_2068_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6753_ (.A1(_2019_),
    .A2(_2031_),
    .ZN(_2069_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6754_ (.A1(_2019_),
    .A2(_2031_),
    .ZN(_2070_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6755_ (.A1(_2017_),
    .A2(_2069_),
    .B(_2070_),
    .ZN(_2071_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6756_ (.A1(_4138_),
    .A2(_1973_),
    .ZN(_2072_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6757_ (.A1(_2022_),
    .A2(_2072_),
    .ZN(_2073_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6758_ (.A1(_4076_),
    .A2(_1902_),
    .ZN(_2074_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6759_ (.A1(_2073_),
    .A2(_2074_),
    .Z(_2075_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6760_ (.A1(_2026_),
    .A2(_2029_),
    .ZN(_2076_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6761_ (.A1(_2023_),
    .A2(_2030_),
    .ZN(_2077_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6762_ (.A1(_2076_),
    .A2(_2077_),
    .ZN(_2078_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6763_ (.A1(_2024_),
    .A2(_2027_),
    .ZN(_2079_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6764_ (.A1(\as2650.r0[3] ),
    .A2(_4089_),
    .ZN(_2080_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6765_ (.A1(_1989_),
    .A2(_2080_),
    .ZN(_2081_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6766_ (.A1(_2079_),
    .A2(_2028_),
    .B(_2081_),
    .ZN(_2082_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6767_ (.A1(\as2650.r0[4] ),
    .A2(_1857_),
    .ZN(_2083_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6768_ (.A1(_2080_),
    .A2(_2083_),
    .ZN(_2084_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6769_ (.A1(_1968_),
    .A2(_1860_),
    .ZN(_2085_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6770_ (.A1(_2084_),
    .A2(_2085_),
    .ZN(_2086_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6771_ (.A1(_2082_),
    .A2(_2086_),
    .Z(_2087_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6772_ (.A1(_2012_),
    .A2(_2087_),
    .Z(_2088_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6773_ (.A1(_2078_),
    .A2(_2088_),
    .Z(_2089_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6774_ (.A1(_2075_),
    .A2(_2089_),
    .Z(_2090_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6775_ (.A1(_2071_),
    .A2(_2090_),
    .Z(_2091_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6776_ (.A1(_2068_),
    .A2(_2091_),
    .ZN(_2092_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6777_ (.A1(_2065_),
    .A2(_2092_),
    .ZN(_2093_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6778_ (.A1(_2063_),
    .A2(_2093_),
    .Z(_2094_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6779_ (.A1(\as2650.r123_2[2][1] ),
    .A2(_1856_),
    .B1(_2094_),
    .B2(_2038_),
    .ZN(_2095_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6780_ (.A1(_1832_),
    .A2(_2061_),
    .B(_2095_),
    .ZN(_0116_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6781_ (.I(_1850_),
    .Z(_2096_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6782_ (.I(_1833_),
    .Z(_2097_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6783_ (.I(_1806_),
    .Z(_2098_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6784_ (.I(_1821_),
    .Z(_2099_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6785_ (.I(_1817_),
    .Z(_2100_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6786_ (.A1(_0882_),
    .A2(_2049_),
    .ZN(_2101_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6787_ (.I(_2046_),
    .Z(_2102_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6788_ (.A1(_4214_),
    .A2(_1814_),
    .B(_2101_),
    .C(_2102_),
    .ZN(_2103_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6789_ (.A1(_4134_),
    .A2(_2048_),
    .B(_2100_),
    .C(_2103_),
    .ZN(_2104_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6790_ (.A1(_0674_),
    .A2(_2045_),
    .B(_2099_),
    .C(_2104_),
    .ZN(_2105_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6791_ (.A1(_0877_),
    .A2(_2042_),
    .B(_1835_),
    .C(_2105_),
    .ZN(_2106_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6792_ (.A1(_0875_),
    .A2(_2098_),
    .B(_2106_),
    .ZN(_2107_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6793_ (.A1(_2097_),
    .A2(_2107_),
    .ZN(_2108_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6794_ (.A1(_0896_),
    .A2(_1826_),
    .ZN(_2109_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6795_ (.A1(_2057_),
    .A2(_2108_),
    .A3(_2109_),
    .ZN(_2110_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6796_ (.A1(_0866_),
    .A2(_2096_),
    .B(_2110_),
    .ZN(_2111_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6797_ (.I(_1855_),
    .Z(_2112_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6798_ (.A1(_2065_),
    .A2(_2092_),
    .Z(_2113_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6799_ (.A1(_2063_),
    .A2(_2093_),
    .B(_2113_),
    .ZN(_2114_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6800_ (.A1(_2071_),
    .A2(_2090_),
    .Z(_2115_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6801_ (.A1(_2068_),
    .A2(_2091_),
    .B(_2115_),
    .ZN(_2116_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6802_ (.A1(_1186_),
    .A2(_2005_),
    .A3(_2073_),
    .ZN(_2117_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _6803_ (.A1(_1954_),
    .A2(_2021_),
    .A3(_2072_),
    .B(_2117_),
    .ZN(_2118_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6804_ (.I(_2088_),
    .ZN(_2119_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6805_ (.A1(_2078_),
    .A2(_2119_),
    .ZN(_2120_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6806_ (.A1(_2075_),
    .A2(_2089_),
    .B(_2120_),
    .ZN(_2121_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6807_ (.A1(_0918_),
    .A2(_2003_),
    .ZN(_2122_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6808_ (.A1(_4100_),
    .A2(_1915_),
    .A3(_2087_),
    .ZN(_2123_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6809_ (.A1(_2082_),
    .A2(_2086_),
    .B(_2123_),
    .ZN(_2124_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6810_ (.A1(_2080_),
    .A2(_2083_),
    .ZN(_2125_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6811_ (.A1(_2084_),
    .A2(_2085_),
    .ZN(_2126_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6812_ (.A1(_2125_),
    .A2(_2126_),
    .ZN(_2127_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6813_ (.A1(\as2650.r0[5] ),
    .A2(_4089_),
    .ZN(_2128_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6814_ (.A1(_2083_),
    .A2(_2128_),
    .ZN(_2129_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6815_ (.A1(_1968_),
    .A2(_1858_),
    .B1(_4090_),
    .B2(\as2650.r0[4] ),
    .ZN(_2130_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6816_ (.A1(_2129_),
    .A2(_2130_),
    .Z(_2131_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6817_ (.A1(_4098_),
    .A2(_1861_),
    .ZN(_2132_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6818_ (.A1(_2131_),
    .A2(_2132_),
    .ZN(_2133_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6819_ (.A1(_2127_),
    .A2(_2133_),
    .Z(_2134_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6820_ (.A1(_2021_),
    .A2(_2134_),
    .ZN(_2135_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6821_ (.A1(_2124_),
    .A2(_2135_),
    .ZN(_2136_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6822_ (.A1(_2122_),
    .A2(_2136_),
    .Z(_2137_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6823_ (.A1(_2121_),
    .A2(_2137_),
    .Z(_2138_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6824_ (.A1(_2118_),
    .A2(_2138_),
    .ZN(_2139_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6825_ (.A1(_2116_),
    .A2(_2139_),
    .Z(_2140_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6826_ (.A1(_2114_),
    .A2(_2140_),
    .Z(_2141_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6827_ (.I(_2037_),
    .Z(_2142_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6828_ (.A1(\as2650.r123_2[2][2] ),
    .A2(_2112_),
    .B1(_2141_),
    .B2(_2142_),
    .ZN(_2143_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6829_ (.A1(_1832_),
    .A2(_2111_),
    .B(_2143_),
    .ZN(_0117_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6830_ (.I(_0951_),
    .Z(_2144_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6831_ (.A1(_0953_),
    .A2(_1813_),
    .ZN(_2145_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6832_ (.A1(_4212_),
    .A2(_1837_),
    .B(_2145_),
    .C(_2047_),
    .ZN(_2146_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6833_ (.A1(_2144_),
    .A2(_2102_),
    .B(_1818_),
    .C(_2146_),
    .ZN(_2147_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6834_ (.A1(_0950_),
    .A2(_2100_),
    .B(_1836_),
    .C(_2147_),
    .ZN(_2148_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6835_ (.A1(_0949_),
    .A2(_2044_),
    .B(_2148_),
    .ZN(_2149_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6836_ (.A1(_2043_),
    .A2(_2149_),
    .ZN(_2150_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6837_ (.A1(_0962_),
    .A2(_2041_),
    .B(_1834_),
    .C(_2150_),
    .ZN(_2151_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6838_ (.A1(_0948_),
    .A2(_2040_),
    .B(_2151_),
    .C(_2057_),
    .ZN(_2152_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6839_ (.A1(_0940_),
    .A2(_2096_),
    .B(_2152_),
    .ZN(_2153_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6840_ (.A1(_2121_),
    .A2(_2137_),
    .ZN(_2154_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6841_ (.A1(_2118_),
    .A2(_2138_),
    .ZN(_2155_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6842_ (.I(_2003_),
    .Z(_2156_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6843_ (.A1(_0988_),
    .A2(_2156_),
    .ZN(_2157_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6844_ (.A1(_4099_),
    .A2(_1864_),
    .ZN(_2158_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6845_ (.I(_2158_),
    .ZN(_2159_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6846_ (.A1(_4075_),
    .A2(_1865_),
    .Z(_2160_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _6847_ (.A1(_2128_),
    .A2(_2159_),
    .A3(_2160_),
    .Z(_2161_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6848_ (.A1(_2131_),
    .A2(_2132_),
    .ZN(_2162_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6849_ (.A1(_2129_),
    .A2(_2162_),
    .ZN(_2163_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6850_ (.A1(_2161_),
    .A2(_2163_),
    .Z(_2164_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6851_ (.A1(_1186_),
    .A2(_1915_),
    .A3(_2134_),
    .ZN(_2165_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6852_ (.A1(_2127_),
    .A2(_2133_),
    .B(_2165_),
    .ZN(_2166_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6853_ (.A1(_2164_),
    .A2(_2166_),
    .Z(_2167_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6854_ (.A1(_2157_),
    .A2(_2167_),
    .ZN(_2168_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6855_ (.A1(_2124_),
    .A2(_2135_),
    .ZN(_2169_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6856_ (.A1(_2122_),
    .A2(_2136_),
    .B(_2169_),
    .ZN(_2170_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6857_ (.A1(_2168_),
    .A2(_2170_),
    .ZN(_2171_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6858_ (.A1(_2154_),
    .A2(_2155_),
    .B(_2171_),
    .ZN(_2172_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _6859_ (.A1(_2154_),
    .A2(_2155_),
    .A3(_2171_),
    .Z(_2173_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6860_ (.A1(_2172_),
    .A2(_2173_),
    .ZN(_2174_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6861_ (.A1(_2116_),
    .A2(_2139_),
    .ZN(_2175_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6862_ (.A1(_2114_),
    .A2(_2140_),
    .B(_2175_),
    .ZN(_2176_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6863_ (.A1(_2174_),
    .A2(_2176_),
    .ZN(_2177_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6864_ (.A1(\as2650.r123_2[2][3] ),
    .A2(_2112_),
    .B1(_2177_),
    .B2(_2142_),
    .ZN(_2178_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6865_ (.A1(_1832_),
    .A2(_2153_),
    .B(_2178_),
    .ZN(_0118_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6866_ (.A1(_2168_),
    .A2(_2170_),
    .ZN(_2179_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6867_ (.A1(_1087_),
    .A2(_2156_),
    .ZN(_2180_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6868_ (.A1(_2161_),
    .A2(_2163_),
    .Z(_2181_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6869_ (.A1(_4099_),
    .A2(_4091_),
    .ZN(_2182_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6870_ (.A1(_4076_),
    .A2(_1864_),
    .ZN(_2183_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6871_ (.A1(_2182_),
    .A2(_2183_),
    .Z(_2184_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6872_ (.A1(_2128_),
    .A2(_2158_),
    .ZN(_2185_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6873_ (.A1(_2128_),
    .A2(_2158_),
    .ZN(_2186_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6874_ (.A1(_2185_),
    .A2(_2160_),
    .B(_2186_),
    .ZN(_2187_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6875_ (.A1(_2184_),
    .A2(_2187_),
    .Z(_2188_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6876_ (.A1(_2181_),
    .A2(_2188_),
    .ZN(_2189_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6877_ (.A1(_2180_),
    .A2(_2189_),
    .Z(_2190_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6878_ (.A1(_2164_),
    .A2(_2166_),
    .ZN(_2191_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6879_ (.A1(_1017_),
    .A2(_2156_),
    .A3(_2167_),
    .ZN(_2192_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6880_ (.A1(_2191_),
    .A2(_2192_),
    .ZN(_2193_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6881_ (.A1(_2190_),
    .A2(_2193_),
    .ZN(_2194_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6882_ (.A1(_2179_),
    .A2(_2194_),
    .ZN(_2195_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _6883_ (.A1(_2114_),
    .A2(_2140_),
    .B(_2172_),
    .C(_2175_),
    .ZN(_2196_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6884_ (.A1(_2173_),
    .A2(_2196_),
    .ZN(_2197_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6885_ (.A1(_2195_),
    .A2(_2197_),
    .Z(_2198_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6886_ (.A1(_1009_),
    .A2(_2059_),
    .ZN(_2199_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6887_ (.A1(_1022_),
    .A2(_2049_),
    .ZN(_2200_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6888_ (.A1(_4198_),
    .A2(_1814_),
    .B(_2200_),
    .C(_2102_),
    .ZN(_2201_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6889_ (.A1(_4202_),
    .A2(_2048_),
    .B(_2100_),
    .C(_2201_),
    .ZN(_2202_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6890_ (.A1(_0880_),
    .A2(_2045_),
    .B(_2099_),
    .C(_2202_),
    .ZN(_2203_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6891_ (.A1(_1017_),
    .A2(_2042_),
    .B(_2203_),
    .ZN(_2204_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6892_ (.A1(_2098_),
    .A2(_2204_),
    .ZN(_2205_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6893_ (.A1(_1035_),
    .A2(_2041_),
    .B(_2097_),
    .C(_2205_),
    .ZN(_2206_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6894_ (.A1(_1015_),
    .A2(_1826_),
    .ZN(_2207_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6895_ (.A1(_2057_),
    .A2(_2206_),
    .A3(_2207_),
    .ZN(_2208_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6896_ (.A1(_2199_),
    .A2(_2208_),
    .ZN(_2209_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6897_ (.A1(_1830_),
    .A2(_2209_),
    .ZN(_2210_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6898_ (.A1(\as2650.r123_2[2][4] ),
    .A2(_1856_),
    .B(_2210_),
    .ZN(_2211_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _6899_ (.A1(_0740_),
    .A2(_1812_),
    .A3(_2198_),
    .B(_2211_),
    .ZN(_0119_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6900_ (.I(_1104_),
    .ZN(_2212_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6901_ (.A1(_1094_),
    .A2(_2049_),
    .ZN(_2213_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6902_ (.A1(_4204_),
    .A2(_1837_),
    .B(_2213_),
    .C(_2047_),
    .ZN(_2214_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6903_ (.A1(_1668_),
    .A2(_2048_),
    .B(_1818_),
    .C(_2214_),
    .ZN(_2215_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6904_ (.A1(_1099_),
    .A2(_2045_),
    .B(_2099_),
    .C(_2215_),
    .ZN(_2216_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6905_ (.A1(_1087_),
    .A2(_2044_),
    .B(_1835_),
    .C(_2216_),
    .ZN(_2217_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6906_ (.A1(_2212_),
    .A2(_2098_),
    .B(_2217_),
    .ZN(_2218_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6907_ (.A1(_2097_),
    .A2(_2218_),
    .ZN(_2219_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6908_ (.A1(_1086_),
    .A2(_1826_),
    .B(_2059_),
    .ZN(_2220_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6909_ (.A1(_1078_),
    .A2(_2059_),
    .B1(_2219_),
    .B2(_2220_),
    .ZN(_2221_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6910_ (.I(_2221_),
    .ZN(_2222_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6911_ (.A1(_2190_),
    .A2(_2193_),
    .ZN(_2223_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6912_ (.A1(_2179_),
    .A2(_2194_),
    .Z(_2224_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _6913_ (.A1(_2173_),
    .A2(_2195_),
    .A3(_2196_),
    .B(_2224_),
    .ZN(_2225_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6914_ (.I(_2187_),
    .ZN(_2226_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6915_ (.A1(_2184_),
    .A2(_2226_),
    .ZN(_2227_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6916_ (.A1(_1186_),
    .A2(_4092_),
    .A3(_2158_),
    .ZN(_2228_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6917_ (.A1(_2227_),
    .A2(_2228_),
    .ZN(_2229_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6918_ (.I(_2156_),
    .Z(_2230_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6919_ (.A1(_1120_),
    .A2(_2230_),
    .ZN(_2231_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6920_ (.A1(_2229_),
    .A2(_2231_),
    .Z(_2232_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _6921_ (.A1(_2161_),
    .A2(_2163_),
    .A3(_2188_),
    .B1(_2189_),
    .B2(_2180_),
    .ZN(_2233_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6922_ (.A1(_2232_),
    .A2(_2233_),
    .Z(_2234_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6923_ (.I(_2234_),
    .ZN(_2235_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _6924_ (.A1(_2223_),
    .A2(_2225_),
    .A3(_2235_),
    .Z(_2236_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6925_ (.A1(\as2650.r123_2[2][5] ),
    .A2(_2112_),
    .B1(_2236_),
    .B2(_2142_),
    .ZN(_2237_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6926_ (.A1(_1831_),
    .A2(_2222_),
    .B(_2237_),
    .ZN(_0120_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6927_ (.I(_1138_),
    .ZN(_2238_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6928_ (.A1(_1144_),
    .A2(_1840_),
    .ZN(_2239_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6929_ (.A1(_1659_),
    .A2(_1814_),
    .B(_1811_),
    .ZN(_2240_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6930_ (.A1(_4081_),
    .A2(_1811_),
    .B1(_2239_),
    .B2(_2240_),
    .ZN(_2241_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6931_ (.A1(_4202_),
    .A2(_1842_),
    .ZN(_2242_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6932_ (.A1(_1842_),
    .A2(_2241_),
    .B(_2242_),
    .C(_2099_),
    .ZN(_2243_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6933_ (.A1(_1121_),
    .A2(_2042_),
    .B(_2043_),
    .C(_2243_),
    .ZN(_2244_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6934_ (.A1(_2238_),
    .A2(_2041_),
    .B(_2097_),
    .C(_2244_),
    .ZN(_2245_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6935_ (.A1(_1154_),
    .A2(_2040_),
    .B(_2245_),
    .ZN(_2246_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6936_ (.I0(_1177_),
    .I1(_2246_),
    .S(_2096_),
    .Z(_2247_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6937_ (.A1(_2223_),
    .A2(_2235_),
    .ZN(_2248_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6938_ (.A1(_2223_),
    .A2(_2235_),
    .ZN(_2249_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6939_ (.A1(_2225_),
    .A2(_2248_),
    .B(_2249_),
    .ZN(_2250_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6940_ (.A1(_2232_),
    .A2(_2233_),
    .ZN(_2251_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6941_ (.A1(_2227_),
    .A2(_2228_),
    .ZN(_2252_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6942_ (.A1(_2229_),
    .A2(_2231_),
    .ZN(_2253_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6943_ (.A1(_2252_),
    .A2(_2253_),
    .ZN(_2254_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _6944_ (.A1(_1187_),
    .A2(_2230_),
    .A3(_4092_),
    .A4(_2159_),
    .ZN(_2255_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6945_ (.A1(_1187_),
    .A2(_2230_),
    .ZN(_2256_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6946_ (.A1(_2182_),
    .A2(_2183_),
    .B(_2256_),
    .ZN(_2257_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6947_ (.A1(_2255_),
    .A2(_2257_),
    .ZN(_2258_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6948_ (.A1(_2254_),
    .A2(_2258_),
    .ZN(_2259_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6949_ (.A1(_2251_),
    .A2(_2259_),
    .ZN(_2260_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6950_ (.A1(_2250_),
    .A2(_2260_),
    .Z(_2261_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6951_ (.A1(\as2650.r123_2[2][6] ),
    .A2(_2112_),
    .B1(_2261_),
    .B2(_2142_),
    .ZN(_2262_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6952_ (.A1(_1831_),
    .A2(_2247_),
    .B(_2262_),
    .ZN(_0121_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6953_ (.I(_1214_),
    .Z(_2263_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6954_ (.A1(_2263_),
    .A2(_1840_),
    .ZN(_2264_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6955_ (.A1(_1217_),
    .A2(_1840_),
    .B(_2264_),
    .C(_1810_),
    .ZN(_2265_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6956_ (.A1(_1213_),
    .A2(_2102_),
    .B(_1817_),
    .ZN(_2266_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _6957_ (.A1(_1089_),
    .A2(_2100_),
    .B1(_2265_),
    .B2(_2266_),
    .C(_1836_),
    .ZN(_2267_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6958_ (.A1(_1210_),
    .A2(_2044_),
    .B(_2267_),
    .ZN(_2268_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6959_ (.A1(_2043_),
    .A2(_2268_),
    .ZN(_2269_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6960_ (.A1(_1228_),
    .A2(_2098_),
    .B(_1834_),
    .C(_2269_),
    .ZN(_2270_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6961_ (.A1(_1234_),
    .A2(_2040_),
    .B(_2270_),
    .C(_1850_),
    .ZN(_2271_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6962_ (.A1(_1209_),
    .A2(_2096_),
    .B(_2271_),
    .ZN(_2272_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6963_ (.A1(_2251_),
    .A2(_2259_),
    .ZN(_2273_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6964_ (.A1(_2254_),
    .A2(_2258_),
    .B(_2255_),
    .ZN(_2274_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6965_ (.A1(_2273_),
    .A2(_2274_),
    .ZN(_2275_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6966_ (.A1(_2250_),
    .A2(_2260_),
    .B(_2275_),
    .ZN(_2276_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6967_ (.A1(_2038_),
    .A2(_2276_),
    .ZN(_2277_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6968_ (.A1(\as2650.r123_2[2][7] ),
    .A2(_1856_),
    .ZN(_2278_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6969_ (.A1(_1831_),
    .A2(_2272_),
    .B(_2277_),
    .C(_2278_),
    .ZN(_0122_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6970_ (.I(_1283_),
    .Z(_2279_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6971_ (.I(_1366_),
    .Z(_2280_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6972_ (.A1(_2280_),
    .A2(_0711_),
    .A3(_1270_),
    .ZN(_2281_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6973_ (.I(_2281_),
    .Z(_2282_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6974_ (.I(_2281_),
    .Z(_2283_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6975_ (.A1(\as2650.stack[5][0] ),
    .A2(_2283_),
    .ZN(_2284_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6976_ (.A1(_2279_),
    .A2(_2282_),
    .B(_2284_),
    .ZN(_0123_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6977_ (.I(_1289_),
    .Z(_2285_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6978_ (.A1(\as2650.stack[5][1] ),
    .A2(_2283_),
    .ZN(_2286_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6979_ (.A1(_2285_),
    .A2(_2282_),
    .B(_2286_),
    .ZN(_0124_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6980_ (.I(_1293_),
    .Z(_2287_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6981_ (.A1(\as2650.stack[5][2] ),
    .A2(_2283_),
    .ZN(_2288_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6982_ (.A1(_2287_),
    .A2(_2282_),
    .B(_2288_),
    .ZN(_0125_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6983_ (.I(_1299_),
    .Z(_2289_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6984_ (.A1(\as2650.stack[5][3] ),
    .A2(_2283_),
    .ZN(_2290_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6985_ (.A1(_2289_),
    .A2(_2282_),
    .B(_2290_),
    .ZN(_0126_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6986_ (.I(_1308_),
    .Z(_2291_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6987_ (.I(_2281_),
    .Z(_2292_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6988_ (.I(_2281_),
    .Z(_2293_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6989_ (.A1(\as2650.stack[5][4] ),
    .A2(_2293_),
    .ZN(_2294_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6990_ (.A1(_2291_),
    .A2(_2292_),
    .B(_2294_),
    .ZN(_0127_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6991_ (.I(_1316_),
    .Z(_2295_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6992_ (.A1(\as2650.stack[5][5] ),
    .A2(_2293_),
    .ZN(_2296_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6993_ (.A1(_2295_),
    .A2(_2292_),
    .B(_2296_),
    .ZN(_0128_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6994_ (.I(_1324_),
    .Z(_2297_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6995_ (.A1(\as2650.stack[5][6] ),
    .A2(_2293_),
    .ZN(_2298_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6996_ (.A1(_2297_),
    .A2(_2292_),
    .B(_2298_),
    .ZN(_0129_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6997_ (.I(_1330_),
    .Z(_2299_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6998_ (.A1(\as2650.stack[5][7] ),
    .A2(_2293_),
    .ZN(_2300_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6999_ (.A1(_2299_),
    .A2(_2292_),
    .B(_2300_),
    .ZN(_0130_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7000_ (.A1(_1633_),
    .A2(_1829_),
    .ZN(_2301_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7001_ (.I(_2301_),
    .Z(_2302_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7002_ (.A1(_1633_),
    .A2(_1829_),
    .B(_1854_),
    .C(_0322_),
    .ZN(_2303_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7003_ (.I(_2303_),
    .Z(_2304_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7004_ (.A1(_2038_),
    .A2(_1924_),
    .B1(_2304_),
    .B2(\as2650.r123_2[1][0] ),
    .ZN(_2305_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7005_ (.A1(_1852_),
    .A2(_2302_),
    .B(_2305_),
    .ZN(_0131_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7006_ (.I(_2303_),
    .Z(_2306_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7007_ (.A1(_0778_),
    .A2(_1923_),
    .ZN(_2307_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7008_ (.A1(_1897_),
    .A2(_2307_),
    .ZN(_2308_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7009_ (.A1(_1927_),
    .A2(_2308_),
    .Z(_2309_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7010_ (.I(_2037_),
    .Z(_2310_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7011_ (.A1(\as2650.r123_2[1][1] ),
    .A2(_2306_),
    .B1(_2309_),
    .B2(_2310_),
    .ZN(_2311_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7012_ (.A1(_2061_),
    .A2(_2302_),
    .B(_2311_),
    .ZN(_0132_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7013_ (.A1(_1928_),
    .A2(_1930_),
    .Z(_2312_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7014_ (.A1(\as2650.r123_2[1][2] ),
    .A2(_2306_),
    .B1(_2312_),
    .B2(_2310_),
    .ZN(_2313_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7015_ (.A1(_2111_),
    .A2(_2302_),
    .B(_2313_),
    .ZN(_0133_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7016_ (.A1(_1932_),
    .A2(_1933_),
    .Z(_2314_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7017_ (.A1(\as2650.r123_2[1][3] ),
    .A2(_2306_),
    .B1(_2314_),
    .B2(_2310_),
    .ZN(_2315_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7018_ (.A1(_2153_),
    .A2(_2302_),
    .B(_2315_),
    .ZN(_0134_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7019_ (.I(_2301_),
    .Z(_2316_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7020_ (.A1(_1921_),
    .A2(_1934_),
    .Z(_2317_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7021_ (.A1(\as2650.r123_2[1][4] ),
    .A2(_2306_),
    .B1(_2317_),
    .B2(_2310_),
    .ZN(_2318_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7022_ (.A1(_2209_),
    .A2(_2316_),
    .B(_2318_),
    .ZN(_0135_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _7023_ (.A1(_1920_),
    .A2(_1935_),
    .A3(_1936_),
    .Z(_2319_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7024_ (.A1(_1937_),
    .A2(_2319_),
    .ZN(_2320_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7025_ (.I(_1854_),
    .Z(_2321_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7026_ (.A1(\as2650.r123_2[1][5] ),
    .A2(_2304_),
    .B1(_2320_),
    .B2(_2321_),
    .ZN(_2322_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7027_ (.A1(_2222_),
    .A2(_2316_),
    .B(_2322_),
    .ZN(_0136_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _7028_ (.A1(_1909_),
    .A2(_1937_),
    .A3(_1960_),
    .Z(_2323_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7029_ (.A1(_1961_),
    .A2(_2323_),
    .Z(_2324_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7030_ (.A1(\as2650.r123_2[1][6] ),
    .A2(_2304_),
    .B1(_2324_),
    .B2(_2321_),
    .ZN(_2325_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7031_ (.A1(_2247_),
    .A2(_2316_),
    .B(_2325_),
    .ZN(_0137_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7032_ (.A1(_1961_),
    .A2(_1996_),
    .Z(_2326_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7033_ (.A1(\as2650.r123_2[1][7] ),
    .A2(_2304_),
    .B1(_2326_),
    .B2(_2321_),
    .ZN(_2327_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7034_ (.A1(_2272_),
    .A2(_2316_),
    .B(_2327_),
    .ZN(_0138_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7035_ (.I(_1708_),
    .Z(_2328_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7036_ (.I(_2328_),
    .Z(_2329_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7037_ (.I(_0562_),
    .Z(_2330_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7038_ (.I(_2330_),
    .Z(_2331_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7039_ (.A1(_0443_),
    .A2(_4275_),
    .ZN(_2332_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7040_ (.A1(_2331_),
    .A2(_1764_),
    .A3(_2332_),
    .ZN(_2333_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7041_ (.I(_4447_),
    .Z(_2334_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7042_ (.I(_2334_),
    .Z(_2335_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7043_ (.I(_1245_),
    .Z(_2336_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _7044_ (.A1(_4360_),
    .A2(_2335_),
    .A3(_2336_),
    .A4(_0389_),
    .ZN(_2337_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _7045_ (.A1(_4046_),
    .A2(_4270_),
    .A3(_1244_),
    .ZN(_2338_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7046_ (.A1(_2337_),
    .A2(_2338_),
    .B(_4401_),
    .ZN(_2339_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7047_ (.A1(_1587_),
    .A2(_1519_),
    .ZN(_2340_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7048_ (.A1(_1518_),
    .A2(_2340_),
    .B(_0434_),
    .C(_1514_),
    .ZN(_2341_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7049_ (.A1(_4256_),
    .A2(_4287_),
    .A3(_0552_),
    .ZN(_2342_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _7050_ (.A1(_0353_),
    .A2(_4341_),
    .A3(_0562_),
    .ZN(_2343_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7051_ (.A1(_1518_),
    .A2(_1520_),
    .Z(_2344_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7052_ (.A1(_4265_),
    .A2(_4337_),
    .Z(_2345_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7053_ (.A1(_0329_),
    .A2(_2345_),
    .B(_0323_),
    .ZN(_2346_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7054_ (.A1(_0404_),
    .A2(_2346_),
    .ZN(_2347_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7055_ (.A1(_2344_),
    .A2(_2347_),
    .ZN(_2348_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7056_ (.A1(_4323_),
    .A2(_0516_),
    .ZN(_2349_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _7057_ (.A1(_2342_),
    .A2(_2343_),
    .A3(_2348_),
    .A4(_2349_),
    .ZN(_2350_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7058_ (.A1(_2341_),
    .A2(_2350_),
    .ZN(_2351_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7059_ (.I(_0359_),
    .Z(_2352_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7060_ (.A1(_2352_),
    .A2(_4346_),
    .ZN(_2353_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7061_ (.I(_2353_),
    .Z(_2354_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7062_ (.I(_4448_),
    .Z(_2355_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7063_ (.A1(_1473_),
    .A2(_2355_),
    .ZN(_2356_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7064_ (.A1(_1488_),
    .A2(_0361_),
    .B1(_2354_),
    .B2(_2356_),
    .ZN(_2357_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _7065_ (.A1(_2333_),
    .A2(_2339_),
    .A3(_2351_),
    .A4(_2357_),
    .ZN(_2358_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7066_ (.I(_2358_),
    .Z(_2359_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7067_ (.I(_2359_),
    .Z(_2360_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7068_ (.I(\as2650.addr_buff[0] ),
    .Z(_2361_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7069_ (.I(_2361_),
    .Z(_2362_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7070_ (.I(_2358_),
    .Z(_2363_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7071_ (.A1(_2362_),
    .A2(_2363_),
    .ZN(_2364_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7072_ (.A1(_2329_),
    .A2(_2360_),
    .B(_2364_),
    .ZN(_0139_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7073_ (.I(_1713_),
    .Z(_2365_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7074_ (.I(\as2650.addr_buff[1] ),
    .Z(_2366_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7075_ (.I(_2358_),
    .Z(_2367_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7076_ (.A1(_2366_),
    .A2(_2367_),
    .ZN(_2368_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7077_ (.A1(_2365_),
    .A2(_2360_),
    .B(_2368_),
    .ZN(_0140_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7078_ (.I(_1718_),
    .Z(_2369_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7079_ (.I(\as2650.addr_buff[2] ),
    .Z(_2370_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7080_ (.I(_2370_),
    .Z(_2371_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7081_ (.A1(_2371_),
    .A2(_2367_),
    .ZN(_2372_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7082_ (.A1(_2369_),
    .A2(_2360_),
    .B(_2372_),
    .ZN(_0141_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7083_ (.I(_1710_),
    .Z(_2373_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7084_ (.I(\as2650.addr_buff[3] ),
    .Z(_2374_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7085_ (.A1(_2374_),
    .A2(_2367_),
    .ZN(_2375_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7086_ (.A1(_2373_),
    .A2(_2360_),
    .B(_2375_),
    .ZN(_0142_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7087_ (.I(_1672_),
    .Z(_2376_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7088_ (.I(_2376_),
    .Z(_2377_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7089_ (.I(\as2650.addr_buff[4] ),
    .Z(_2378_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7090_ (.I0(_2377_),
    .I1(_2378_),
    .S(_2359_),
    .Z(_2379_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7091_ (.I(_2379_),
    .Z(_0143_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7092_ (.I(_0533_),
    .Z(_2380_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7093_ (.A1(_2380_),
    .A2(_2367_),
    .ZN(_2381_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7094_ (.A1(_1502_),
    .A2(_2363_),
    .B(_2381_),
    .ZN(_0144_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7095_ (.I(_0532_),
    .Z(_2382_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7096_ (.A1(_2382_),
    .A2(_2359_),
    .ZN(_2383_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7097_ (.A1(_1659_),
    .A2(_2363_),
    .B(_2383_),
    .ZN(_0145_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7098_ (.I(_1216_),
    .Z(_2384_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7099_ (.I(_2384_),
    .Z(_2385_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7100_ (.A1(_4432_),
    .A2(_2359_),
    .ZN(_2386_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7101_ (.A1(_2385_),
    .A2(_2363_),
    .B(_2386_),
    .ZN(_0146_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7102_ (.A1(_0706_),
    .A2(_0702_),
    .ZN(_2387_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7103_ (.I(_2387_),
    .Z(_2388_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7104_ (.I(_2388_),
    .Z(_2389_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _7105_ (.A1(_1243_),
    .A2(_2389_),
    .A3(_1782_),
    .ZN(_2390_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7106_ (.I(_2390_),
    .Z(_2391_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7107_ (.I(_2391_),
    .Z(_2392_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7108_ (.I(_2391_),
    .Z(_2393_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7109_ (.A1(\as2650.stack[4][8] ),
    .A2(_2393_),
    .ZN(_2394_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7110_ (.A1(_1781_),
    .A2(_2392_),
    .B(_2394_),
    .ZN(_0147_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7111_ (.I(_2390_),
    .Z(_2395_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7112_ (.A1(\as2650.stack[4][9] ),
    .A2(_2395_),
    .ZN(_2396_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7113_ (.A1(_1789_),
    .A2(_2392_),
    .B(_2396_),
    .ZN(_0148_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7114_ (.A1(\as2650.stack[4][10] ),
    .A2(_2395_),
    .ZN(_2397_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7115_ (.A1(_1792_),
    .A2(_2392_),
    .B(_2397_),
    .ZN(_0149_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7116_ (.A1(\as2650.stack[4][11] ),
    .A2(_2395_),
    .ZN(_2398_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7117_ (.A1(_1794_),
    .A2(_2392_),
    .B(_2398_),
    .ZN(_0150_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7118_ (.A1(\as2650.stack[4][12] ),
    .A2(_2395_),
    .ZN(_2399_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7119_ (.A1(_1796_),
    .A2(_2393_),
    .B(_2399_),
    .ZN(_0151_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7120_ (.A1(\as2650.stack[4][13] ),
    .A2(_2391_),
    .ZN(_2400_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7121_ (.A1(_1798_),
    .A2(_2393_),
    .B(_2400_),
    .ZN(_0152_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7122_ (.A1(\as2650.stack[4][14] ),
    .A2(_2391_),
    .ZN(_2401_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7123_ (.A1(_1800_),
    .A2(_2393_),
    .B(_2401_),
    .ZN(_0153_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7124_ (.I(_0573_),
    .Z(_2402_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7125_ (.A1(_1131_),
    .A2(_1828_),
    .ZN(_2403_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _7126_ (.A1(_2402_),
    .A2(_1815_),
    .B(_2403_),
    .C(_4343_),
    .ZN(_2404_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7127_ (.I(_2404_),
    .Z(_2405_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7128_ (.I(_2403_),
    .Z(_2406_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7129_ (.I(_0737_),
    .Z(_2407_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7130_ (.A1(_2407_),
    .A2(_0815_),
    .A3(_1808_),
    .ZN(_2408_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7131_ (.I(_2408_),
    .Z(_2409_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7132_ (.I(_0732_),
    .Z(_2410_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7133_ (.A1(_2410_),
    .A2(_1815_),
    .ZN(_2411_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _7134_ (.A1(_0663_),
    .A2(_2411_),
    .Z(_2412_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7135_ (.A1(_0730_),
    .A2(_2409_),
    .B(_2412_),
    .ZN(_2413_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7136_ (.A1(_2402_),
    .A2(_1815_),
    .ZN(_2414_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7137_ (.A1(_1854_),
    .A2(_2414_),
    .ZN(_2415_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7138_ (.I(_2404_),
    .Z(_2416_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _7139_ (.A1(_1852_),
    .A2(_2406_),
    .B1(_2413_),
    .B2(_2415_),
    .C(_2416_),
    .ZN(_2417_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7140_ (.A1(\as2650.r123_2[0][0] ),
    .A2(_2405_),
    .B(_2417_),
    .ZN(_2418_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7141_ (.I(_2418_),
    .ZN(_0154_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7142_ (.I(_2403_),
    .Z(_2419_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7143_ (.I(_2404_),
    .Z(_2420_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7144_ (.I(_1853_),
    .Z(_2421_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7145_ (.I(_2414_),
    .Z(_2422_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7146_ (.I(_2411_),
    .Z(_2423_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _7147_ (.A1(_0832_),
    .A2(_2409_),
    .Z(_2424_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _7148_ (.A1(_2421_),
    .A2(_2422_),
    .B1(_2423_),
    .B2(_1540_),
    .C(_2424_),
    .ZN(_2425_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7149_ (.A1(_2061_),
    .A2(_2419_),
    .B(_2420_),
    .C(_2425_),
    .ZN(_2426_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7150_ (.A1(\as2650.r123_2[0][1] ),
    .A2(_2405_),
    .B(_2426_),
    .ZN(_2427_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7151_ (.I(_2427_),
    .ZN(_0155_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7152_ (.I(_2408_),
    .Z(_2428_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _7153_ (.A1(_0908_),
    .A2(_2428_),
    .Z(_2429_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _7154_ (.A1(_2421_),
    .A2(_2422_),
    .B1(_2423_),
    .B2(_1545_),
    .C(_2429_),
    .ZN(_2430_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7155_ (.A1(_2111_),
    .A2(_2419_),
    .B(_2420_),
    .C(_2430_),
    .ZN(_2431_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7156_ (.A1(\as2650.r123_2[0][2] ),
    .A2(_2405_),
    .B(_2431_),
    .ZN(_2432_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7157_ (.I(_2432_),
    .ZN(_0156_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _7158_ (.A1(_0978_),
    .A2(_2428_),
    .Z(_2433_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _7159_ (.A1(_2421_),
    .A2(_2422_),
    .B1(_2423_),
    .B2(_0969_),
    .C(_2433_),
    .ZN(_2434_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7160_ (.A1(_2153_),
    .A2(_2419_),
    .B(_2420_),
    .C(_2434_),
    .ZN(_2435_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7161_ (.A1(\as2650.r123_2[0][3] ),
    .A2(_2405_),
    .B(_2435_),
    .ZN(_2436_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7162_ (.I(_2436_),
    .ZN(_0157_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7163_ (.I(_2404_),
    .Z(_2437_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _7164_ (.A1(_1049_),
    .A2(_2428_),
    .Z(_2438_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _7165_ (.A1(_2421_),
    .A2(_2414_),
    .B1(_2411_),
    .B2(_1303_),
    .C(_2438_),
    .ZN(_2439_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7166_ (.A1(_2209_),
    .A2(_2406_),
    .B(_2416_),
    .C(_2439_),
    .ZN(_2440_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7167_ (.A1(\as2650.r123_2[0][4] ),
    .A2(_2437_),
    .B(_2440_),
    .ZN(_2441_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7168_ (.I(_2441_),
    .ZN(_0158_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _7169_ (.A1(_1114_),
    .A2(_2428_),
    .Z(_2442_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _7170_ (.A1(_2037_),
    .A2(_2414_),
    .B1(_2411_),
    .B2(_1312_),
    .C(_2442_),
    .ZN(_2443_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7171_ (.A1(_2222_),
    .A2(_2406_),
    .B(_2416_),
    .C(_2443_),
    .ZN(_2444_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7172_ (.A1(\as2650.r123_2[0][5] ),
    .A2(_2437_),
    .B(_2444_),
    .ZN(_2445_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7173_ (.I(_2445_),
    .ZN(_0159_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _7174_ (.A1(\as2650.r123_2[0][6] ),
    .A2(_2420_),
    .Z(_2446_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _7175_ (.A1(_1128_),
    .A2(_2409_),
    .Z(_2447_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _7176_ (.A1(_2321_),
    .A2(_2422_),
    .B1(_2423_),
    .B2(_1319_),
    .C(_2447_),
    .ZN(_2448_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7177_ (.A1(_2247_),
    .A2(_2419_),
    .B(_2437_),
    .C(_2448_),
    .ZN(_2449_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7178_ (.A1(_2446_),
    .A2(_2449_),
    .Z(_2450_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7179_ (.I(_2450_),
    .Z(_0160_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7180_ (.A1(_1211_),
    .A2(_2409_),
    .ZN(_2451_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _7181_ (.A1(_2272_),
    .A2(_2406_),
    .B1(_2415_),
    .B2(_2451_),
    .C(_2416_),
    .ZN(_2452_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7182_ (.A1(\as2650.r123_2[0][7] ),
    .A2(_2437_),
    .B(_2452_),
    .ZN(_2453_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7183_ (.I(_2453_),
    .ZN(_0161_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7184_ (.A1(_0706_),
    .A2(\as2650.psu[1] ),
    .ZN(_2454_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7185_ (.I(_2454_),
    .Z(_2455_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7186_ (.I(_2455_),
    .Z(_2456_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _7187_ (.A1(_1366_),
    .A2(_2456_),
    .A3(_1367_),
    .ZN(_2457_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7188_ (.I(_2457_),
    .Z(_2458_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7189_ (.I(_2458_),
    .Z(_2459_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7190_ (.I(_2458_),
    .Z(_2460_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7191_ (.A1(\as2650.stack[2][8] ),
    .A2(_2460_),
    .ZN(_2461_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7192_ (.A1(_2459_),
    .A2(_1386_),
    .B(_2461_),
    .ZN(_0162_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7193_ (.I(_2457_),
    .Z(_2462_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7194_ (.A1(\as2650.stack[2][9] ),
    .A2(_2462_),
    .ZN(_2463_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7195_ (.A1(_2459_),
    .A2(_1396_),
    .B(_2463_),
    .ZN(_0163_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7196_ (.A1(\as2650.stack[2][10] ),
    .A2(_2462_),
    .ZN(_2464_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7197_ (.A1(_2459_),
    .A2(_1404_),
    .B(_2464_),
    .ZN(_0164_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7198_ (.A1(\as2650.stack[2][11] ),
    .A2(_2462_),
    .ZN(_2465_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7199_ (.A1(_2459_),
    .A2(_1414_),
    .B(_2465_),
    .ZN(_0165_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7200_ (.A1(\as2650.stack[2][12] ),
    .A2(_2462_),
    .ZN(_2466_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7201_ (.A1(_2460_),
    .A2(_1420_),
    .B(_2466_),
    .ZN(_0166_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7202_ (.A1(\as2650.stack[2][13] ),
    .A2(_2458_),
    .ZN(_2467_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7203_ (.A1(_2460_),
    .A2(_1427_),
    .B(_2467_),
    .ZN(_0167_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7204_ (.A1(\as2650.stack[2][14] ),
    .A2(_2458_),
    .ZN(_2468_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7205_ (.A1(_2460_),
    .A2(_1434_),
    .B(_2468_),
    .ZN(_0168_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7206_ (.A1(_1526_),
    .A2(_2343_),
    .ZN(_2469_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7207_ (.A1(_0451_),
    .A2(_2340_),
    .ZN(_2470_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7208_ (.I(_0812_),
    .Z(_2471_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7209_ (.I(_2471_),
    .Z(_2472_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7210_ (.I(_2472_),
    .Z(_2473_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _7211_ (.A1(_2473_),
    .A2(_4353_),
    .A3(_0291_),
    .ZN(_2474_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _7212_ (.A1(_1517_),
    .A2(_2469_),
    .A3(_2470_),
    .A4(_2474_),
    .ZN(_2475_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7213_ (.A1(_4354_),
    .A2(_0387_),
    .B(_0307_),
    .ZN(_2476_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7214_ (.A1(net25),
    .A2(_2475_),
    .ZN(_2477_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7215_ (.A1(_2475_),
    .A2(_2476_),
    .B(_2477_),
    .C(_1568_),
    .ZN(_0169_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7216_ (.I(_1246_),
    .Z(_2478_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _7217_ (.A1(_0341_),
    .A2(_1468_),
    .A3(_0481_),
    .ZN(_2479_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7218_ (.A1(_2478_),
    .A2(_2479_),
    .ZN(_2480_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _7219_ (.A1(_0465_),
    .A2(_4051_),
    .A3(_2480_),
    .ZN(_2481_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7220_ (.I(_1686_),
    .Z(_2482_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7221_ (.A1(net23),
    .A2(_2481_),
    .B(_2482_),
    .ZN(_2483_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7222_ (.A1(_4392_),
    .A2(_2481_),
    .B(_2483_),
    .ZN(_0170_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7223_ (.I(net24),
    .ZN(_2484_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7224_ (.A1(_1635_),
    .A2(_2479_),
    .B(_0339_),
    .ZN(_2485_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7225_ (.I(_1253_),
    .Z(_2486_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _7226_ (.A1(_4353_),
    .A2(_2486_),
    .A3(_1629_),
    .Z(_2487_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _7227_ (.A1(_4323_),
    .A2(_1253_),
    .ZN(_2488_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _7228_ (.A1(_4353_),
    .A2(_1477_),
    .A3(_0291_),
    .A4(_2488_),
    .ZN(_2489_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _7229_ (.A1(_0465_),
    .A2(_2485_),
    .A3(_2487_),
    .A4(_2489_),
    .ZN(_2490_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7230_ (.A1(_4051_),
    .A2(_0340_),
    .B(_2490_),
    .ZN(_2491_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7231_ (.A1(_2484_),
    .A2(_2490_),
    .B(_2491_),
    .C(_1689_),
    .ZN(_0171_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7232_ (.A1(_4348_),
    .A2(_4284_),
    .ZN(_2492_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7233_ (.A1(_0550_),
    .A2(_0561_),
    .ZN(_2493_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _7234_ (.A1(_4387_),
    .A2(_2493_),
    .ZN(_2494_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7235_ (.A1(_2492_),
    .A2(_2494_),
    .ZN(_2495_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _7236_ (.A1(_0317_),
    .A2(_4340_),
    .A3(_2495_),
    .ZN(_2496_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7237_ (.I(_1512_),
    .Z(_2497_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7238_ (.I(_1247_),
    .Z(_2498_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7239_ (.A1(_2497_),
    .A2(_2498_),
    .ZN(_2499_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7240_ (.A1(_0471_),
    .A2(_1266_),
    .ZN(_2500_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7241_ (.A1(_4237_),
    .A2(_1278_),
    .ZN(_2501_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7242_ (.I(_2501_),
    .ZN(_2502_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7243_ (.A1(_0739_),
    .A2(_1279_),
    .B1(_2338_),
    .B2(_2502_),
    .ZN(_2503_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _7244_ (.A1(_0353_),
    .A2(_4346_),
    .B(_0556_),
    .C(_1513_),
    .ZN(_2504_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7245_ (.A1(_4441_),
    .A2(_1481_),
    .A3(_1459_),
    .ZN(_2505_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7246_ (.A1(_4322_),
    .A2(_4329_),
    .A3(_1253_),
    .ZN(_2506_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _7247_ (.A1(_2503_),
    .A2(_2504_),
    .A3(_2505_),
    .A4(_2506_),
    .Z(_2507_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7248_ (.A1(_4308_),
    .A2(_1481_),
    .ZN(_2508_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7249_ (.A1(_1649_),
    .A2(_1278_),
    .ZN(_2509_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7250_ (.A1(_0483_),
    .A2(_1278_),
    .ZN(_2510_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _7251_ (.A1(_1643_),
    .A2(_1266_),
    .B1(_2509_),
    .B2(_0475_),
    .C(_2510_),
    .ZN(_2511_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _7252_ (.A1(_0310_),
    .A2(_2494_),
    .B(_1749_),
    .C(_4290_),
    .ZN(_2512_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _7253_ (.A1(_4283_),
    .A2(_4348_),
    .A3(_0556_),
    .A4(_1520_),
    .ZN(_2513_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7254_ (.A1(_2512_),
    .A2(_2513_),
    .ZN(_2514_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7255_ (.A1(_4298_),
    .A2(_0491_),
    .B(_0486_),
    .C(_0501_),
    .ZN(_2515_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7256_ (.A1(_1279_),
    .A2(_2515_),
    .ZN(_2516_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7257_ (.A1(_0731_),
    .A2(_2509_),
    .B(_2516_),
    .ZN(_2517_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7258_ (.I(_2493_),
    .Z(_2518_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7259_ (.A1(_4405_),
    .A2(_2518_),
    .ZN(_2519_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _7260_ (.A1(_4276_),
    .A2(_2332_),
    .A3(_2519_),
    .Z(_2520_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _7261_ (.A1(_2511_),
    .A2(_2514_),
    .A3(_2517_),
    .A4(_2520_),
    .ZN(_2521_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _7262_ (.A1(_2480_),
    .A2(_2507_),
    .A3(_2508_),
    .A4(_2521_),
    .ZN(_2522_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _7263_ (.A1(_2496_),
    .A2(_2499_),
    .A3(_2500_),
    .A4(_2522_),
    .ZN(_2523_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7264_ (.I(_2523_),
    .Z(_2524_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7265_ (.I(_2524_),
    .Z(_2525_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7266_ (.I(_2525_),
    .Z(_2526_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7267_ (.I(_1277_),
    .Z(_2527_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7268_ (.A1(_4401_),
    .A2(_2478_),
    .ZN(_2528_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7269_ (.A1(_1252_),
    .A2(_2528_),
    .ZN(_2529_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7270_ (.I(_2529_),
    .Z(_2530_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7271_ (.I(_0376_),
    .Z(_2531_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7272_ (.A1(_0813_),
    .A2(_4439_),
    .ZN(_2532_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7273_ (.A1(_2531_),
    .A2(_2532_),
    .ZN(_2533_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7274_ (.I(_2533_),
    .Z(_2534_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7275_ (.A1(_2527_),
    .A2(_0321_),
    .ZN(_2535_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7276_ (.I(_1215_),
    .Z(_2536_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7277_ (.I(_2536_),
    .Z(_2537_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7278_ (.I(_2537_),
    .Z(_2538_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7279_ (.A1(_1276_),
    .A2(_2328_),
    .Z(_2539_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7280_ (.I(net29),
    .Z(_2540_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7281_ (.I(_2540_),
    .Z(_2541_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7282_ (.I(_2384_),
    .Z(_2542_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7283_ (.A1(_2541_),
    .A2(_2542_),
    .ZN(_2543_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7284_ (.A1(_4441_),
    .A2(_0397_),
    .ZN(_2544_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7285_ (.A1(_2471_),
    .A2(_2544_),
    .ZN(_2545_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7286_ (.I(_2545_),
    .Z(_2546_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7287_ (.A1(_2538_),
    .A2(_2539_),
    .B(_2543_),
    .C(_2546_),
    .ZN(_2547_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7288_ (.I(_4442_),
    .Z(_2548_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _7289_ (.A1(_1479_),
    .A2(_0358_),
    .A3(_2548_),
    .ZN(_2549_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7290_ (.I(_4430_),
    .Z(_2550_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7291_ (.I(_2550_),
    .Z(_2551_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7292_ (.I(_4434_),
    .Z(_2552_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7293_ (.I(_2552_),
    .Z(_2553_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7294_ (.I(_4411_),
    .Z(_2554_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7295_ (.I(_2554_),
    .Z(_2555_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7296_ (.A1(_2555_),
    .A2(_2328_),
    .ZN(_2556_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7297_ (.A1(_2540_),
    .A2(_2551_),
    .B(_2553_),
    .C(_2556_),
    .ZN(_2557_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7298_ (.A1(_2541_),
    .A2(_4437_),
    .B(_2549_),
    .C(_2557_),
    .ZN(_2558_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7299_ (.A1(_2547_),
    .A2(_2558_),
    .B(_4242_),
    .ZN(_2559_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7300_ (.A1(_4430_),
    .A2(_1531_),
    .ZN(_2560_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7301_ (.I(_2560_),
    .Z(_2561_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7302_ (.I(_2561_),
    .Z(_2562_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7303_ (.A1(_1752_),
    .A2(_0660_),
    .A3(_2562_),
    .ZN(_2563_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7304_ (.I(_2560_),
    .Z(_2564_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7305_ (.A1(_0660_),
    .A2(_2564_),
    .ZN(_2565_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7306_ (.I(_0326_),
    .Z(_2566_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7307_ (.A1(_2329_),
    .A2(_2565_),
    .B(_2566_),
    .C(_0419_),
    .ZN(_2567_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7308_ (.I(_0641_),
    .Z(_2568_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _7309_ (.A1(_1708_),
    .A2(_0650_),
    .Z(_2569_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7310_ (.A1(_2568_),
    .A2(_2569_),
    .ZN(_2570_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7311_ (.I(_4339_),
    .Z(_2571_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7312_ (.A1(_2568_),
    .A2(_0651_),
    .B(_2328_),
    .ZN(_2572_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7313_ (.A1(_4336_),
    .A2(_2571_),
    .A3(_2572_),
    .ZN(_2573_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7314_ (.A1(_4048_),
    .A2(_1509_),
    .ZN(_2574_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7315_ (.A1(_4409_),
    .A2(_2539_),
    .B(_2574_),
    .ZN(_2575_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _7316_ (.A1(_2541_),
    .A2(_2347_),
    .B1(_2570_),
    .B2(_2573_),
    .C(_2575_),
    .ZN(_2576_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7317_ (.A1(_2563_),
    .A2(_2567_),
    .B(_2576_),
    .ZN(_2577_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7318_ (.A1(_2534_),
    .A2(_2535_),
    .B(_2559_),
    .C(_2577_),
    .ZN(_2578_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7319_ (.A1(_2527_),
    .A2(_2530_),
    .B1(_2578_),
    .B2(_0458_),
    .ZN(_2579_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7320_ (.A1(_2541_),
    .A2(_2525_),
    .ZN(_2580_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7321_ (.A1(_2526_),
    .A2(_2579_),
    .B(_2580_),
    .C(_1568_),
    .ZN(_0172_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7322_ (.I(_2524_),
    .Z(_2581_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7323_ (.I(\as2650.pc[1] ),
    .Z(_2582_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7324_ (.I(_2529_),
    .Z(_2583_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7325_ (.I(net3),
    .Z(_2584_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7326_ (.I(_2584_),
    .Z(_2585_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7327_ (.I(_2585_),
    .Z(_2586_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7328_ (.I(_2586_),
    .Z(_2587_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7329_ (.A1(_1274_),
    .A2(net7),
    .ZN(_2588_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7330_ (.A1(\as2650.pc[1] ),
    .A2(net8),
    .ZN(_2589_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7331_ (.A1(_2588_),
    .A2(_2589_),
    .Z(_2590_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7332_ (.A1(_2587_),
    .A2(_2590_),
    .ZN(_2591_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7333_ (.I(net30),
    .Z(_2592_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7334_ (.A1(_2592_),
    .A2(_2538_),
    .ZN(_2593_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7335_ (.A1(_2546_),
    .A2(_2591_),
    .A3(_2593_),
    .ZN(_2594_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7336_ (.A1(_4324_),
    .A2(_4313_),
    .ZN(_2595_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7337_ (.I(_2595_),
    .Z(_2596_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7338_ (.I(_2596_),
    .Z(_2597_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7339_ (.A1(_1499_),
    .A2(_2597_),
    .B(_1288_),
    .ZN(_2598_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7340_ (.A1(_2592_),
    .A2(_2540_),
    .ZN(_2599_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7341_ (.I(_2552_),
    .Z(_2600_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7342_ (.I(_2554_),
    .Z(_2601_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7343_ (.A1(_2601_),
    .A2(_2365_),
    .ZN(_2602_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7344_ (.A1(_2592_),
    .A2(_2551_),
    .B(_2600_),
    .C(_2602_),
    .ZN(_2603_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7345_ (.A1(_4437_),
    .A2(_2599_),
    .B(_2603_),
    .C(_2549_),
    .ZN(_2604_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7346_ (.A1(_2594_),
    .A2(_2598_),
    .A3(_2604_),
    .ZN(_2605_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7347_ (.I(_4276_),
    .Z(_2606_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7348_ (.I(_0404_),
    .Z(_2607_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7349_ (.A1(_0785_),
    .A2(_0801_),
    .Z(_2608_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7350_ (.A1(_0676_),
    .A2(_0659_),
    .B(_2608_),
    .ZN(_2609_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7351_ (.A1(_0675_),
    .A2(_0659_),
    .A3(_2608_),
    .ZN(_2610_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7352_ (.A1(_2560_),
    .A2(_2610_),
    .ZN(_2611_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7353_ (.I(_2345_),
    .Z(_2612_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _7354_ (.A1(_1713_),
    .A2(_2561_),
    .B1(_2609_),
    .B2(_2611_),
    .C(_2612_),
    .ZN(_2613_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7355_ (.I(_0542_),
    .Z(_2614_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7356_ (.A1(_1712_),
    .A2(_0806_),
    .Z(_2615_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7357_ (.A1(_2569_),
    .A2(_2615_),
    .Z(_2616_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7358_ (.A1(_2614_),
    .A2(_2616_),
    .ZN(_2617_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7359_ (.A1(_1713_),
    .A2(_2614_),
    .B(_2617_),
    .C(_4339_),
    .ZN(_2618_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7360_ (.A1(_2613_),
    .A2(_2618_),
    .ZN(_2619_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7361_ (.I(_2346_),
    .Z(_2620_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7362_ (.A1(_0324_),
    .A2(_2619_),
    .B1(_2599_),
    .B2(_2620_),
    .ZN(_2621_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7363_ (.A1(\as2650.pc[0] ),
    .A2(net7),
    .ZN(_2622_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _7364_ (.A1(_2622_),
    .A2(_2589_),
    .Z(_2623_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7365_ (.A1(_2622_),
    .A2(_2589_),
    .B(_0405_),
    .ZN(_2624_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _7366_ (.A1(_2607_),
    .A2(_2621_),
    .B1(_2623_),
    .B2(_2624_),
    .C(_2574_),
    .ZN(_2625_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7367_ (.A1(_1288_),
    .A2(_0380_),
    .B1(_2605_),
    .B2(_2606_),
    .C(_2625_),
    .ZN(_2626_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7368_ (.A1(_2582_),
    .A2(_2583_),
    .B1(_2626_),
    .B2(_0458_),
    .ZN(_2627_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7369_ (.A1(_2592_),
    .A2(_2525_),
    .ZN(_2628_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7370_ (.I(_1507_),
    .Z(_2629_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7371_ (.A1(_2581_),
    .A2(_2627_),
    .B(_2628_),
    .C(_2629_),
    .ZN(_0173_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7372_ (.I(net31),
    .Z(_2630_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7373_ (.A1(net30),
    .A2(_2540_),
    .ZN(_2631_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7374_ (.A1(_2630_),
    .A2(_2631_),
    .Z(_2632_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7375_ (.A1(\as2650.pc[2] ),
    .A2(net9),
    .Z(_2633_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7376_ (.I(_2633_),
    .Z(_2634_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7377_ (.A1(\as2650.pc[1] ),
    .A2(_0784_),
    .ZN(_2635_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7378_ (.A1(_2635_),
    .A2(_2623_),
    .ZN(_2636_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7379_ (.A1(_2634_),
    .A2(_2636_),
    .Z(_2637_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7380_ (.A1(_0417_),
    .A2(_2637_),
    .ZN(_2638_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7381_ (.I(_0883_),
    .Z(_2639_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7382_ (.A1(_0785_),
    .A2(_0806_),
    .ZN(_2640_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _7383_ (.A1(_2569_),
    .A2(_2615_),
    .B(_2640_),
    .ZN(_2641_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _7384_ (.A1(_0893_),
    .A2(_0895_),
    .B(_1717_),
    .ZN(_2642_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7385_ (.A1(_0883_),
    .A2(_0896_),
    .ZN(_2643_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7386_ (.A1(_2642_),
    .A2(_2643_),
    .ZN(_2644_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7387_ (.A1(_2641_),
    .A2(_2644_),
    .B(_0641_),
    .ZN(_2645_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7388_ (.A1(_2641_),
    .A2(_2644_),
    .B(_2645_),
    .ZN(_2646_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7389_ (.A1(_2639_),
    .A2(_2614_),
    .B(_2646_),
    .C(_2571_),
    .ZN(_2647_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7390_ (.A1(_0786_),
    .A2(_0802_),
    .ZN(_2648_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7391_ (.A1(_2648_),
    .A2(_2610_),
    .ZN(_2649_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _7392_ (.A1(_0882_),
    .A2(_0874_),
    .ZN(_2650_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7393_ (.A1(_1718_),
    .A2(_0875_),
    .ZN(_2651_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _7394_ (.A1(_2649_),
    .A2(_2650_),
    .A3(_2651_),
    .ZN(_2652_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7395_ (.A1(_2650_),
    .A2(_2651_),
    .B(_2649_),
    .ZN(_2653_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7396_ (.A1(_2561_),
    .A2(_2653_),
    .ZN(_2654_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _7397_ (.A1(_2639_),
    .A2(_2561_),
    .B1(_2652_),
    .B2(_2654_),
    .C(_2612_),
    .ZN(_2655_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7398_ (.A1(_2647_),
    .A2(_2655_),
    .ZN(_2656_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7399_ (.A1(_4336_),
    .A2(_2656_),
    .ZN(_2657_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7400_ (.A1(_2347_),
    .A2(_2632_),
    .B(_2638_),
    .C(_2657_),
    .ZN(_2658_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7401_ (.A1(_2588_),
    .A2(_2589_),
    .B(_2635_),
    .ZN(_2659_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7402_ (.A1(_2634_),
    .A2(_2659_),
    .ZN(_2660_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7403_ (.A1(_2630_),
    .A2(_0412_),
    .B(_2546_),
    .ZN(_2661_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7404_ (.A1(_1694_),
    .A2(_2660_),
    .B(_2661_),
    .ZN(_2662_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7405_ (.I(\as2650.pc[2] ),
    .Z(_2663_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7406_ (.I(_2663_),
    .Z(_2664_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7407_ (.A1(_2664_),
    .A2(_0305_),
    .A3(_2533_),
    .ZN(_2665_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7408_ (.I(_2335_),
    .Z(_2666_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7409_ (.A1(_2551_),
    .A2(_2639_),
    .ZN(_2667_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7410_ (.A1(_2630_),
    .A2(_0461_),
    .B(_2355_),
    .ZN(_2668_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7411_ (.A1(_2666_),
    .A2(_2632_),
    .B1(_2667_),
    .B2(_2668_),
    .C(_1259_),
    .ZN(_2669_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7412_ (.A1(_1764_),
    .A2(_2669_),
    .ZN(_2670_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7413_ (.A1(_2665_),
    .A2(_2670_),
    .ZN(_2671_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7414_ (.A1(_1588_),
    .A2(_2658_),
    .B1(_2662_),
    .B2(_4276_),
    .C(_2671_),
    .ZN(_2672_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7415_ (.I(_0338_),
    .Z(_2673_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _7416_ (.A1(_1292_),
    .A2(_2583_),
    .B1(_2672_),
    .B2(_2673_),
    .C(_2525_),
    .ZN(_2674_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7417_ (.I(_2523_),
    .Z(_2675_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _7418_ (.A1(_2630_),
    .A2(_2675_),
    .Z(_2676_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _7419_ (.A1(_1689_),
    .A2(_2674_),
    .A3(_2676_),
    .Z(_2677_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7420_ (.I(_2677_),
    .Z(_0174_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7421_ (.I(_0324_),
    .Z(_2678_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _7422_ (.A1(_0944_),
    .A2(_0947_),
    .ZN(_2679_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7423_ (.A1(_1710_),
    .A2(_2679_),
    .Z(_2680_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _7424_ (.A1(_1717_),
    .A2(_0893_),
    .A3(_0895_),
    .ZN(_2681_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7425_ (.A1(_2641_),
    .A2(_2642_),
    .B(_2681_),
    .ZN(_2682_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7426_ (.A1(_2680_),
    .A2(_2682_),
    .B(_2614_),
    .ZN(_2683_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7427_ (.A1(_2680_),
    .A2(_2682_),
    .B(_2683_),
    .ZN(_2684_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7428_ (.I(_0542_),
    .Z(_2685_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7429_ (.I(_4339_),
    .Z(_2686_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7430_ (.A1(_2373_),
    .A2(_2685_),
    .B(_2686_),
    .ZN(_2687_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7431_ (.A1(_0881_),
    .A2(_0874_),
    .ZN(_2688_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _7432_ (.A1(_2648_),
    .A2(_2610_),
    .A3(_2688_),
    .Z(_2689_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7433_ (.A1(_2650_),
    .A2(_2689_),
    .ZN(_2690_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _7434_ (.A1(_1679_),
    .A2(_0962_),
    .A3(_2690_),
    .Z(_2691_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7435_ (.A1(_2564_),
    .A2(_2691_),
    .ZN(_2692_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7436_ (.I(_2345_),
    .Z(_2693_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7437_ (.A1(_2373_),
    .A2(_2564_),
    .B(_2692_),
    .C(_2693_),
    .ZN(_2694_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7438_ (.A1(_2684_),
    .A2(_2687_),
    .B(_2694_),
    .ZN(_2695_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7439_ (.A1(net31),
    .A2(net30),
    .A3(net29),
    .ZN(_2696_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7440_ (.A1(net55),
    .A2(_2696_),
    .Z(_2697_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7441_ (.I(_2620_),
    .Z(_2698_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7442_ (.A1(_2678_),
    .A2(_2695_),
    .B1(_2697_),
    .B2(_2698_),
    .C(_4410_),
    .ZN(_2699_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7443_ (.I(_0404_),
    .Z(_2700_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7444_ (.A1(\as2650.pc[3] ),
    .A2(_0952_),
    .ZN(_2701_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7445_ (.A1(_1296_),
    .A2(_1709_),
    .ZN(_2702_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7446_ (.A1(_2701_),
    .A2(_2702_),
    .ZN(_2703_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7447_ (.A1(_1292_),
    .A2(_1717_),
    .ZN(_2704_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7448_ (.A1(_2634_),
    .A2(_2636_),
    .B(_2704_),
    .ZN(_2705_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7449_ (.A1(_2703_),
    .A2(_2705_),
    .Z(_2706_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7450_ (.A1(_0338_),
    .A2(_2574_),
    .ZN(_2707_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7451_ (.A1(_2700_),
    .A2(_2706_),
    .B(_2707_),
    .ZN(_2708_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7452_ (.A1(_2699_),
    .A2(_2708_),
    .ZN(_2709_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7453_ (.I(\as2650.pc[3] ),
    .Z(_2710_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7454_ (.I(net55),
    .ZN(_2711_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7455_ (.I(_0434_),
    .Z(_2712_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7456_ (.A1(_0425_),
    .A2(_0357_),
    .ZN(_2713_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7457_ (.A1(_2712_),
    .A2(_2713_),
    .ZN(_2714_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7458_ (.I(_2585_),
    .Z(_2715_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7459_ (.A1(_2634_),
    .A2(_2659_),
    .B(_2704_),
    .ZN(_2716_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7460_ (.A1(_2703_),
    .A2(_2716_),
    .ZN(_2717_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7461_ (.A1(_2715_),
    .A2(_2717_),
    .ZN(_2718_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7462_ (.A1(_2711_),
    .A2(_2587_),
    .B(_2714_),
    .C(_2718_),
    .ZN(_2719_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7463_ (.I(_4434_),
    .Z(_2720_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7464_ (.I(_2720_),
    .Z(_2721_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7465_ (.I(_2721_),
    .Z(_2722_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7466_ (.I(_4435_),
    .Z(_2723_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7467_ (.A1(_4431_),
    .A2(_1710_),
    .ZN(_2724_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7468_ (.A1(net55),
    .A2(_2601_),
    .B(_2723_),
    .C(_2724_),
    .ZN(_2725_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7469_ (.A1(_2722_),
    .A2(_2697_),
    .B(_2725_),
    .C(_0440_),
    .ZN(_2726_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7470_ (.A1(_2719_),
    .A2(_2726_),
    .ZN(_2727_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7471_ (.I(_2532_),
    .Z(_2728_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7472_ (.I(_2728_),
    .Z(_2729_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7473_ (.A1(_1298_),
    .A2(_2533_),
    .B1(_2727_),
    .B2(_2729_),
    .ZN(_2730_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7474_ (.I(_2528_),
    .Z(_2731_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7475_ (.A1(_2710_),
    .A2(_2529_),
    .B1(_2730_),
    .B2(_2731_),
    .ZN(_2732_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7476_ (.A1(_2709_),
    .A2(_2732_),
    .B(_2675_),
    .ZN(_2733_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7477_ (.A1(net55),
    .A2(_2581_),
    .B(_2733_),
    .ZN(_2734_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7478_ (.A1(_0335_),
    .A2(_2734_),
    .ZN(_0175_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7479_ (.A1(_1304_),
    .A2(net11),
    .Z(_2735_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7480_ (.I(net10),
    .Z(_2736_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7481_ (.A1(_2710_),
    .A2(_2736_),
    .ZN(_2737_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7482_ (.A1(_2701_),
    .A2(_2705_),
    .B(_2737_),
    .ZN(_2738_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7483_ (.A1(_2735_),
    .A2(_2738_),
    .Z(_2739_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7484_ (.I(net33),
    .Z(_2740_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7485_ (.A1(_2711_),
    .A2(_2696_),
    .ZN(_2741_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7486_ (.A1(_2740_),
    .A2(_2741_),
    .Z(_2742_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7487_ (.A1(_0406_),
    .A2(_2698_),
    .A3(_2742_),
    .ZN(_2743_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7488_ (.I(_0639_),
    .Z(_2744_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7489_ (.I(_2568_),
    .Z(_2745_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7490_ (.A1(_2736_),
    .A2(_2679_),
    .ZN(_2746_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _7491_ (.A1(_2736_),
    .A2(_2679_),
    .B1(_2641_),
    .B2(_2642_),
    .C(_2681_),
    .ZN(_2747_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7492_ (.A1(_1019_),
    .A2(_1014_),
    .ZN(_2748_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7493_ (.A1(_2746_),
    .A2(_2747_),
    .B(_2748_),
    .ZN(_2749_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _7494_ (.A1(_2746_),
    .A2(_2748_),
    .A3(_2747_),
    .ZN(_2750_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7495_ (.A1(_2745_),
    .A2(_2750_),
    .ZN(_2751_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7496_ (.A1(_2376_),
    .A2(_2745_),
    .B1(_2749_),
    .B2(_2751_),
    .ZN(_2752_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7497_ (.A1(_2744_),
    .A2(_2752_),
    .ZN(_2753_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7498_ (.A1(_2736_),
    .A2(_0961_),
    .ZN(_2754_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7499_ (.A1(_0953_),
    .A2(_0961_),
    .ZN(_2755_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _7500_ (.A1(_2650_),
    .A2(_2754_),
    .A3(_2689_),
    .B(_2755_),
    .ZN(_2756_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _7501_ (.A1(_1023_),
    .A2(_1035_),
    .A3(_2756_),
    .Z(_2757_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7502_ (.A1(_2562_),
    .A2(_2757_),
    .ZN(_2758_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _7503_ (.A1(_4411_),
    .A2(_1531_),
    .Z(_2759_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7504_ (.I(_2759_),
    .Z(_2760_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7505_ (.A1(_2376_),
    .A2(_2760_),
    .ZN(_2761_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7506_ (.I(_0326_),
    .Z(_2762_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7507_ (.A1(_2758_),
    .A2(_2761_),
    .B(_2762_),
    .ZN(_2763_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7508_ (.A1(_2753_),
    .A2(_2763_),
    .B(_4336_),
    .ZN(_2764_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7509_ (.A1(_0406_),
    .A2(_2739_),
    .B(_2743_),
    .C(_2764_),
    .ZN(_2765_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7510_ (.I(\as2650.pc[4] ),
    .Z(_2766_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7511_ (.I(_2766_),
    .Z(_2767_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7512_ (.I(_0460_),
    .Z(_2768_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7513_ (.A1(_2740_),
    .A2(_2768_),
    .ZN(_2769_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7514_ (.A1(_2555_),
    .A2(_1672_),
    .ZN(_2770_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7515_ (.A1(_2600_),
    .A2(_2769_),
    .A3(_2770_),
    .ZN(_2771_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7516_ (.A1(_2722_),
    .A2(_2742_),
    .B(_2771_),
    .C(_0441_),
    .ZN(_2772_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7517_ (.A1(_2766_),
    .A2(net11),
    .Z(_2773_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7518_ (.A1(_2633_),
    .A2(_2659_),
    .B(_2702_),
    .C(_2704_),
    .ZN(_2774_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _7519_ (.A1(_2701_),
    .A2(_2774_),
    .Z(_2775_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7520_ (.A1(_2773_),
    .A2(_2775_),
    .Z(_2776_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7521_ (.A1(_1693_),
    .A2(_2776_),
    .ZN(_2777_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7522_ (.A1(_2740_),
    .A2(_0393_),
    .B(_2714_),
    .C(_2777_),
    .ZN(_2778_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7523_ (.A1(_2772_),
    .A2(_2778_),
    .ZN(_2779_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7524_ (.A1(_2767_),
    .A2(_2534_),
    .B1(_2779_),
    .B2(_2729_),
    .ZN(_2780_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7525_ (.I(_2528_),
    .Z(_2781_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7526_ (.I(_2781_),
    .Z(_2782_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _7527_ (.A1(_1305_),
    .A2(_2583_),
    .B1(_2780_),
    .B2(_2782_),
    .C(_2675_),
    .ZN(_2783_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7528_ (.A1(_2707_),
    .A2(_2765_),
    .B(_2783_),
    .ZN(_2784_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7529_ (.A1(_2740_),
    .A2(_2581_),
    .B(_1687_),
    .ZN(_2785_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7530_ (.A1(_2784_),
    .A2(_2785_),
    .ZN(_0176_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7531_ (.I(_2524_),
    .Z(_2786_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7532_ (.I(_2786_),
    .Z(_2787_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7533_ (.I(\as2650.pc[5] ),
    .Z(_2788_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7534_ (.I(_2788_),
    .Z(_2789_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7535_ (.A1(_1313_),
    .A2(_1091_),
    .Z(_2790_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7536_ (.A1(_2766_),
    .A2(_1021_),
    .ZN(_2791_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7537_ (.A1(_2773_),
    .A2(_2738_),
    .ZN(_2792_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7538_ (.A1(_2791_),
    .A2(_2792_),
    .ZN(_2793_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7539_ (.A1(_2790_),
    .A2(_2793_),
    .Z(_2794_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7540_ (.I(_0314_),
    .Z(_2795_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7541_ (.A1(_1490_),
    .A2(_2760_),
    .ZN(_2796_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _7542_ (.A1(_1020_),
    .A2(_1034_),
    .Z(_2797_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7543_ (.A1(_1020_),
    .A2(_1034_),
    .Z(_2798_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7544_ (.A1(_2797_),
    .A2(_2756_),
    .B(_2798_),
    .ZN(_2799_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _7545_ (.A1(_1501_),
    .A2(_1104_),
    .A3(_2799_),
    .Z(_2800_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7546_ (.A1(_2562_),
    .A2(_2800_),
    .B(_0326_),
    .ZN(_2801_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7547_ (.A1(_1490_),
    .A2(_2745_),
    .B(_2744_),
    .ZN(_2802_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7548_ (.A1(_1020_),
    .A2(_1015_),
    .ZN(_2803_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _7549_ (.A1(_2746_),
    .A2(_2748_),
    .A3(_2747_),
    .B(_2803_),
    .ZN(_2804_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _7550_ (.A1(_1094_),
    .A2(_1086_),
    .A3(_2804_),
    .Z(_2805_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7551_ (.A1(_2685_),
    .A2(_2805_),
    .ZN(_2806_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7552_ (.A1(_2796_),
    .A2(_2801_),
    .B1(_2802_),
    .B2(_2806_),
    .ZN(_2807_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7553_ (.I(_2346_),
    .Z(_2808_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7554_ (.I(net34),
    .Z(_2809_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7555_ (.A1(net33),
    .A2(_2741_),
    .Z(_2810_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7556_ (.A1(_2809_),
    .A2(_2810_),
    .ZN(_2811_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7557_ (.A1(_2808_),
    .A2(_2811_),
    .ZN(_2812_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7558_ (.A1(_2795_),
    .A2(_2807_),
    .B(_2812_),
    .C(_2607_),
    .ZN(_2813_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7559_ (.I(_1587_),
    .Z(_2814_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7560_ (.A1(_0406_),
    .A2(_2794_),
    .B(_2813_),
    .C(_2814_),
    .ZN(_2815_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7561_ (.I(_2528_),
    .Z(_2816_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7562_ (.A1(_2788_),
    .A2(_1091_),
    .Z(_2817_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7563_ (.A1(_2735_),
    .A2(_2775_),
    .B(_2791_),
    .ZN(_2818_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7564_ (.A1(_2817_),
    .A2(_2818_),
    .Z(_2819_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7565_ (.I0(_2809_),
    .I1(_2819_),
    .S(_2715_),
    .Z(_2820_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7566_ (.I(_2554_),
    .Z(_2821_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7567_ (.A1(_2821_),
    .A2(_1502_),
    .ZN(_2822_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7568_ (.A1(_2809_),
    .A2(_2601_),
    .B(_2723_),
    .C(_2822_),
    .ZN(_2823_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7569_ (.A1(_2722_),
    .A2(_2811_),
    .B(_2823_),
    .C(_0440_),
    .ZN(_2824_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7570_ (.A1(_2544_),
    .A2(_2820_),
    .B(_2824_),
    .ZN(_2825_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7571_ (.A1(_1314_),
    .A2(_2534_),
    .B1(_2825_),
    .B2(_2729_),
    .ZN(_2826_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _7572_ (.A1(_2816_),
    .A2(_2826_),
    .Z(_2827_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _7573_ (.A1(_2789_),
    .A2(_2530_),
    .B1(_2815_),
    .B2(_0458_),
    .C(_2827_),
    .ZN(_2828_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7574_ (.I(_2524_),
    .Z(_2829_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7575_ (.I(_0350_),
    .Z(_2830_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7576_ (.A1(_2809_),
    .A2(_2829_),
    .B(_2830_),
    .ZN(_2831_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7577_ (.A1(_2787_),
    .A2(_2828_),
    .B(_2831_),
    .ZN(_0177_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7578_ (.I(net35),
    .Z(_2832_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7579_ (.A1(_1657_),
    .A2(_1137_),
    .Z(_2833_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7580_ (.A1(_1093_),
    .A2(_1103_),
    .ZN(_2834_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _7581_ (.A1(_1093_),
    .A2(_1103_),
    .B1(_2797_),
    .B2(_2756_),
    .C(_2798_),
    .ZN(_2835_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7582_ (.A1(_2834_),
    .A2(_2835_),
    .ZN(_2836_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7583_ (.A1(_2833_),
    .A2(_2836_),
    .Z(_2837_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7584_ (.A1(_1673_),
    .A2(_2760_),
    .ZN(_2838_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7585_ (.A1(_2760_),
    .A2(_2837_),
    .B(_2838_),
    .C(_2693_),
    .ZN(_2839_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7586_ (.I(_1140_),
    .Z(_2840_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7587_ (.A1(_2840_),
    .A2(_1153_),
    .Z(_2841_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7588_ (.A1(_1093_),
    .A2(_1085_),
    .Z(_2842_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _7589_ (.A1(_1092_),
    .A2(_1085_),
    .Z(_2843_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7590_ (.A1(_2842_),
    .A2(_2804_),
    .B(_2843_),
    .ZN(_2844_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7591_ (.A1(_2841_),
    .A2(_2844_),
    .Z(_2845_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7592_ (.A1(_1673_),
    .A2(_2568_),
    .ZN(_2846_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7593_ (.A1(_2745_),
    .A2(_2845_),
    .B(_2846_),
    .C(_2571_),
    .ZN(_2847_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7594_ (.A1(_2839_),
    .A2(_2847_),
    .B(_0314_),
    .ZN(_2848_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7595_ (.A1(net34),
    .A2(_2810_),
    .ZN(_2849_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7596_ (.A1(_2832_),
    .A2(_2849_),
    .Z(_2850_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7597_ (.A1(_2620_),
    .A2(_2850_),
    .ZN(_2851_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7598_ (.A1(_0405_),
    .A2(_2851_),
    .ZN(_2852_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7599_ (.A1(\as2650.pc[6] ),
    .A2(_1656_),
    .Z(_2853_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7600_ (.I(_2853_),
    .Z(_2854_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7601_ (.A1(_2792_),
    .A2(_2790_),
    .ZN(_2855_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7602_ (.A1(_2766_),
    .A2(net11),
    .B1(_1091_),
    .B2(_2788_),
    .ZN(_2856_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7603_ (.A1(_1313_),
    .A2(_1500_),
    .B(_2856_),
    .ZN(_2857_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7604_ (.A1(_2855_),
    .A2(_2857_),
    .ZN(_2858_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7605_ (.A1(_2854_),
    .A2(_2858_),
    .ZN(_2859_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _7606_ (.A1(_2848_),
    .A2(_2852_),
    .B1(_2859_),
    .B2(_2607_),
    .C(_1588_),
    .ZN(_2860_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7607_ (.I(_4440_),
    .Z(_2861_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7608_ (.A1(_2832_),
    .A2(_0461_),
    .ZN(_2862_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7609_ (.I(_4447_),
    .Z(_2863_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7610_ (.I(_2863_),
    .Z(_2864_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7611_ (.A1(_2601_),
    .A2(_1673_),
    .B(_2864_),
    .ZN(_2865_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7612_ (.A1(_2666_),
    .A2(_2850_),
    .B1(_2862_),
    .B2(_2865_),
    .ZN(_2866_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7613_ (.A1(_2735_),
    .A2(_2775_),
    .ZN(_2867_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7614_ (.A1(_2867_),
    .A2(_2817_),
    .B(_2857_),
    .ZN(_2868_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7615_ (.A1(_2854_),
    .A2(_2868_),
    .ZN(_2869_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7616_ (.A1(_2832_),
    .A2(_2715_),
    .ZN(_2870_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7617_ (.A1(_2587_),
    .A2(_2869_),
    .B(_2870_),
    .ZN(_2871_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7618_ (.A1(_0441_),
    .A2(_2866_),
    .B1(_2871_),
    .B2(_2714_),
    .ZN(_2872_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7619_ (.A1(_1322_),
    .A2(_2533_),
    .B(_0320_),
    .ZN(_2873_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _7620_ (.A1(_4362_),
    .A2(_2861_),
    .A3(_2872_),
    .B(_2873_),
    .ZN(_2874_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7621_ (.A1(_2860_),
    .A2(_2874_),
    .B(_2673_),
    .ZN(_2875_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7622_ (.A1(_1322_),
    .A2(_2583_),
    .ZN(_2876_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7623_ (.A1(_2875_),
    .A2(_2876_),
    .B(_2675_),
    .ZN(_2877_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7624_ (.A1(_2832_),
    .A2(_2581_),
    .B(_2877_),
    .ZN(_2878_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7625_ (.A1(_0335_),
    .A2(_2878_),
    .ZN(_0178_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7626_ (.I(\as2650.pc[7] ),
    .Z(_2879_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7627_ (.I(_2529_),
    .Z(_2880_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7628_ (.A1(_1327_),
    .A2(_1140_),
    .Z(_2881_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7629_ (.A1(_1320_),
    .A2(_1141_),
    .ZN(_2882_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7630_ (.A1(_2854_),
    .A2(_2868_),
    .B(_2882_),
    .ZN(_2883_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7631_ (.A1(_2881_),
    .A2(_2883_),
    .ZN(_2884_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7632_ (.I(net54),
    .ZN(_2885_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7633_ (.I(_2545_),
    .Z(_2886_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7634_ (.A1(_2885_),
    .A2(_0412_),
    .B(_2886_),
    .ZN(_2887_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7635_ (.A1(_0394_),
    .A2(_2884_),
    .B(_2887_),
    .ZN(_2888_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7636_ (.A1(net35),
    .A2(net34),
    .A3(_2810_),
    .ZN(_2889_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7637_ (.A1(net54),
    .A2(_2889_),
    .Z(_2890_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7638_ (.I(_2720_),
    .Z(_2891_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7639_ (.A1(_2550_),
    .A2(_2384_),
    .ZN(_2892_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7640_ (.A1(net54),
    .A2(_2821_),
    .B(_2891_),
    .C(_2892_),
    .ZN(_2893_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7641_ (.A1(_2600_),
    .A2(_2890_),
    .B(_2893_),
    .C(_2331_),
    .ZN(_2894_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7642_ (.A1(_2879_),
    .A2(_0377_),
    .B(_2894_),
    .ZN(_2895_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7643_ (.A1(_4443_),
    .A2(_2895_),
    .ZN(_2896_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7644_ (.A1(_2879_),
    .A2(_2729_),
    .B(_2896_),
    .ZN(_2897_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7645_ (.I(_2840_),
    .Z(_2898_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7646_ (.A1(_2898_),
    .A2(_1154_),
    .ZN(_2899_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _7647_ (.A1(_2842_),
    .A2(_2804_),
    .B(_2843_),
    .C(_2841_),
    .ZN(_2900_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7648_ (.A1(_2899_),
    .A2(_2900_),
    .ZN(_2901_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _7649_ (.A1(_1216_),
    .A2(_1234_),
    .A3(_2901_),
    .Z(_2902_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7650_ (.I(_2536_),
    .Z(_2903_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7651_ (.A1(_2903_),
    .A2(_2685_),
    .B(_2571_),
    .ZN(_2904_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7652_ (.A1(_2685_),
    .A2(_2902_),
    .B(_2904_),
    .ZN(_2905_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7653_ (.A1(_2898_),
    .A2(_1138_),
    .ZN(_2906_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _7654_ (.A1(_2834_),
    .A2(_2833_),
    .A3(_2835_),
    .B(_2906_),
    .ZN(_2907_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _7655_ (.A1(_0391_),
    .A2(_1228_),
    .A3(_2907_),
    .Z(_2908_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7656_ (.A1(_2903_),
    .A2(_2564_),
    .B(_2612_),
    .ZN(_2909_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7657_ (.A1(_2562_),
    .A2(_2908_),
    .B(_2909_),
    .ZN(_2910_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7658_ (.A1(_2905_),
    .A2(_2910_),
    .B(_2678_),
    .ZN(_2911_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7659_ (.A1(_2808_),
    .A2(_2890_),
    .B(_4410_),
    .ZN(_2912_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7660_ (.A1(_2854_),
    .A2(_2858_),
    .B(_2882_),
    .ZN(_2913_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7661_ (.A1(_2881_),
    .A2(_2913_),
    .Z(_2914_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7662_ (.A1(_0405_),
    .A2(_2914_),
    .B(_1587_),
    .ZN(_2915_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7663_ (.A1(_2911_),
    .A2(_2912_),
    .B(_2915_),
    .ZN(_2916_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7664_ (.A1(_2606_),
    .A2(_2888_),
    .B1(_2897_),
    .B2(_0306_),
    .C(_2916_),
    .ZN(_2917_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7665_ (.A1(_2879_),
    .A2(_2880_),
    .B1(_2917_),
    .B2(_0340_),
    .ZN(_2918_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7666_ (.A1(net54),
    .A2(_2829_),
    .B(_2830_),
    .ZN(_2919_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7667_ (.A1(_2787_),
    .A2(_2918_),
    .B(_2919_),
    .ZN(_0179_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _7668_ (.A1(_1215_),
    .A2(_1233_),
    .B(_2899_),
    .C(_2900_),
    .ZN(_2920_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _7669_ (.A1(_2263_),
    .A2(_1233_),
    .B(_0640_),
    .ZN(_2921_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7670_ (.A1(_2920_),
    .A2(_2921_),
    .ZN(_2922_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7671_ (.A1(_2361_),
    .A2(_2922_),
    .Z(_2923_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7672_ (.A1(_0390_),
    .A2(_1227_),
    .Z(_2924_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7673_ (.A1(_2584_),
    .A2(_1227_),
    .ZN(_2925_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _7674_ (.A1(_2759_),
    .A2(_2925_),
    .ZN(_2926_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7675_ (.A1(_2907_),
    .A2(_2924_),
    .B(_2926_),
    .ZN(_2927_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7676_ (.A1(_2361_),
    .A2(_2927_),
    .Z(_2928_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7677_ (.I(_2612_),
    .Z(_2929_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7678_ (.A1(_2686_),
    .A2(_2923_),
    .B1(_2928_),
    .B2(_2929_),
    .ZN(_2930_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7679_ (.I(net37),
    .Z(_2931_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7680_ (.A1(_2885_),
    .A2(_2889_),
    .ZN(_2932_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7681_ (.A1(_2931_),
    .A2(_2932_),
    .ZN(_2933_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7682_ (.A1(_2698_),
    .A2(_2933_),
    .ZN(_2934_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7683_ (.A1(_2795_),
    .A2(_2930_),
    .B(_2934_),
    .C(_2700_),
    .ZN(_2935_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7684_ (.A1(\as2650.pc[8] ),
    .A2(_1140_),
    .Z(_2936_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _7685_ (.A1(_2853_),
    .A2(_2881_),
    .Z(_2937_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7686_ (.A1(\as2650.pc[7] ),
    .A2(_1141_),
    .ZN(_2938_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7687_ (.A1(_2858_),
    .A2(_2937_),
    .B(_2938_),
    .C(_2882_),
    .ZN(_2939_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7688_ (.A1(_2936_),
    .A2(_2939_),
    .ZN(_2940_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7689_ (.A1(_2936_),
    .A2(_2939_),
    .ZN(_2941_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7690_ (.A1(_2607_),
    .A2(_2941_),
    .ZN(_2942_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7691_ (.I(_2574_),
    .Z(_2943_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7692_ (.A1(_2940_),
    .A2(_2942_),
    .B(_2943_),
    .ZN(_2944_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7693_ (.A1(_2931_),
    .A2(_0461_),
    .ZN(_2945_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7694_ (.A1(_2551_),
    .A2(_2362_),
    .B(_2864_),
    .ZN(_2946_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7695_ (.A1(_2666_),
    .A2(_2933_),
    .B1(_2945_),
    .B2(_2946_),
    .ZN(_2947_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7696_ (.A1(_0441_),
    .A2(_2947_),
    .ZN(_2948_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7697_ (.A1(_2853_),
    .A2(_2881_),
    .ZN(_2949_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7698_ (.A1(_2857_),
    .A2(_2949_),
    .ZN(_2950_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7699_ (.A1(_2882_),
    .A2(_2938_),
    .A3(_2950_),
    .ZN(_2951_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _7700_ (.A1(_2735_),
    .A2(_2775_),
    .A3(_2790_),
    .A4(_2937_),
    .ZN(_2952_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7701_ (.A1(_2951_),
    .A2(_2952_),
    .B(_2936_),
    .ZN(_2953_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _7702_ (.A1(_2936_),
    .A2(_2951_),
    .A3(_2952_),
    .Z(_2954_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7703_ (.A1(_2953_),
    .A2(_2954_),
    .ZN(_2955_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7704_ (.A1(_2587_),
    .A2(_2955_),
    .ZN(_2956_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7705_ (.A1(_2931_),
    .A2(_0393_),
    .B(_2714_),
    .C(_2956_),
    .ZN(_2957_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7706_ (.A1(_2948_),
    .A2(_2957_),
    .ZN(_2958_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7707_ (.I(_2728_),
    .Z(_2959_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7708_ (.A1(_1381_),
    .A2(_2534_),
    .B1(_2958_),
    .B2(_2959_),
    .ZN(_2960_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7709_ (.I(_0386_),
    .Z(_2961_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7710_ (.A1(_2935_),
    .A2(_2944_),
    .B1(_2960_),
    .B2(_2961_),
    .ZN(_2962_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7711_ (.A1(_1381_),
    .A2(_2880_),
    .B1(_2962_),
    .B2(_0340_),
    .ZN(_2963_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7712_ (.A1(_2931_),
    .A2(_2829_),
    .B(_2830_),
    .ZN(_2964_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7713_ (.A1(_2787_),
    .A2(_2963_),
    .B(_2964_),
    .ZN(_0180_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7714_ (.I(\as2650.pc[9] ),
    .Z(_2965_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7715_ (.A1(_1389_),
    .A2(_2840_),
    .Z(_2966_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7716_ (.A1(_1378_),
    .A2(_2898_),
    .ZN(_2967_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7717_ (.A1(_2967_),
    .A2(_2940_),
    .ZN(_2968_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7718_ (.A1(_2966_),
    .A2(_2968_),
    .ZN(_2969_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7719_ (.I(\as2650.addr_buff[1] ),
    .ZN(_2970_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7720_ (.I(_2970_),
    .Z(_2971_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7721_ (.I(\as2650.addr_buff[0] ),
    .Z(_2972_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _7722_ (.A1(_2907_),
    .A2(_2924_),
    .B(_2926_),
    .C(_2972_),
    .ZN(_2973_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7723_ (.A1(_2971_),
    .A2(_2973_),
    .Z(_2974_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7724_ (.A1(_2972_),
    .A2(_2920_),
    .A3(_2921_),
    .ZN(_2975_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7725_ (.A1(_2971_),
    .A2(_2975_),
    .Z(_2976_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7726_ (.A1(_2566_),
    .A2(_2974_),
    .B1(_2976_),
    .B2(_2744_),
    .ZN(_2977_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7727_ (.I(net38),
    .Z(_2978_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7728_ (.A1(net37),
    .A2(_2932_),
    .ZN(_2979_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7729_ (.A1(_2978_),
    .A2(_2979_),
    .Z(_2980_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7730_ (.A1(_2678_),
    .A2(_2977_),
    .B1(_2980_),
    .B2(_2808_),
    .C(_0417_),
    .ZN(_2981_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7731_ (.A1(_0418_),
    .A2(_2969_),
    .B(_2981_),
    .ZN(_2982_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7732_ (.A1(_2967_),
    .A2(_2953_),
    .ZN(_2983_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7733_ (.A1(_2966_),
    .A2(_2983_),
    .Z(_2984_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7734_ (.A1(_2903_),
    .A2(_2984_),
    .ZN(_2985_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7735_ (.A1(_2978_),
    .A2(_2542_),
    .B(_2985_),
    .ZN(_2986_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7736_ (.A1(_2550_),
    .A2(_2970_),
    .ZN(_2987_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7737_ (.A1(_2978_),
    .A2(_4431_),
    .B(_2721_),
    .C(_2987_),
    .ZN(_2988_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7738_ (.I(_2330_),
    .Z(_2989_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7739_ (.A1(_2553_),
    .A2(_2980_),
    .B(_2988_),
    .C(_2989_),
    .ZN(_2990_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7740_ (.A1(_2965_),
    .A2(_0377_),
    .B(_2990_),
    .ZN(_2991_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7741_ (.A1(_2886_),
    .A2(_2986_),
    .B1(_2991_),
    .B2(_4406_),
    .ZN(_2992_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7742_ (.I(_4440_),
    .Z(_2993_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7743_ (.A1(_2965_),
    .A2(_2959_),
    .B1(_2992_),
    .B2(_2993_),
    .ZN(_2994_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7744_ (.A1(_2814_),
    .A2(_2982_),
    .B1(_2994_),
    .B2(_2961_),
    .ZN(_2995_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7745_ (.I(_2673_),
    .Z(_2996_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7746_ (.A1(_2965_),
    .A2(_2880_),
    .B1(_2995_),
    .B2(_2996_),
    .ZN(_2997_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7747_ (.A1(_2978_),
    .A2(_2829_),
    .B(_2830_),
    .ZN(_2998_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7748_ (.A1(_2787_),
    .A2(_2997_),
    .B(_2998_),
    .ZN(_0181_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7749_ (.I(\as2650.pc[10] ),
    .Z(_2999_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7750_ (.I(_2999_),
    .Z(_3000_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7751_ (.A1(_2971_),
    .A2(_2973_),
    .ZN(_3001_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _7752_ (.A1(\as2650.addr_buff[0] ),
    .A2(\as2650.addr_buff[1] ),
    .A3(\as2650.addr_buff[2] ),
    .Z(_3002_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _7753_ (.A1(_2907_),
    .A2(_2924_),
    .B(_2926_),
    .C(_3002_),
    .ZN(_3003_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7754_ (.A1(_2371_),
    .A2(_3001_),
    .B(_3003_),
    .ZN(_3004_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7755_ (.A1(_2971_),
    .A2(_2975_),
    .ZN(_3005_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _7756_ (.A1(_2920_),
    .A2(_2921_),
    .A3(_3002_),
    .ZN(_3006_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7757_ (.A1(_2371_),
    .A2(_3005_),
    .B(_3006_),
    .ZN(_3007_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7758_ (.A1(_2929_),
    .A2(_3004_),
    .B1(_3007_),
    .B2(_2686_),
    .ZN(_3008_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7759_ (.I(net39),
    .Z(_3009_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7760_ (.A1(net38),
    .A2(net37),
    .A3(_2932_),
    .ZN(_3010_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7761_ (.A1(_3009_),
    .A2(_3010_),
    .Z(_3011_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7762_ (.A1(_2698_),
    .A2(_3011_),
    .ZN(_3012_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7763_ (.A1(_2795_),
    .A2(_3008_),
    .B(_3012_),
    .C(_2700_),
    .ZN(_3013_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7764_ (.A1(_1399_),
    .A2(_1141_),
    .Z(_3014_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7765_ (.I(_3014_),
    .Z(_3015_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7766_ (.A1(\as2650.pc[9] ),
    .A2(_1378_),
    .B(_2840_),
    .ZN(_3016_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7767_ (.I(_3016_),
    .ZN(_3017_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7768_ (.A1(_2940_),
    .A2(_2966_),
    .ZN(_3018_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7769_ (.A1(_3017_),
    .A2(_3018_),
    .ZN(_3019_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7770_ (.A1(_3015_),
    .A2(_3019_),
    .Z(_3020_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7771_ (.A1(_0418_),
    .A2(_3020_),
    .B(_2943_),
    .ZN(_3021_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7772_ (.A1(_2953_),
    .A2(_2966_),
    .ZN(_3022_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7773_ (.A1(_3017_),
    .A2(_3022_),
    .ZN(_3023_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7774_ (.A1(_3015_),
    .A2(_3023_),
    .ZN(_3024_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7775_ (.A1(_3009_),
    .A2(_0393_),
    .B(_2546_),
    .C(_0423_),
    .ZN(_3025_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7776_ (.A1(_1694_),
    .A2(_3024_),
    .B(_3025_),
    .ZN(_3026_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7777_ (.I(_2863_),
    .Z(_3027_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7778_ (.A1(_2555_),
    .A2(_2370_),
    .ZN(_3028_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7779_ (.A1(_3009_),
    .A2(_2768_),
    .B(_2335_),
    .ZN(_3029_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7780_ (.A1(_3027_),
    .A2(_3011_),
    .B1(_3028_),
    .B2(_3029_),
    .ZN(_3030_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7781_ (.A1(_3000_),
    .A2(_2597_),
    .B1(_2331_),
    .B2(_3030_),
    .ZN(_3031_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7782_ (.I(_2336_),
    .Z(_3032_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7783_ (.I(_3032_),
    .Z(_3033_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _7784_ (.A1(_1400_),
    .A2(_2728_),
    .B1(_3031_),
    .B2(_3033_),
    .C(_0305_),
    .ZN(_3034_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7785_ (.A1(_3026_),
    .A2(_3034_),
    .ZN(_3035_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7786_ (.A1(_3013_),
    .A2(_3021_),
    .B(_3035_),
    .ZN(_3036_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7787_ (.A1(_3000_),
    .A2(_2880_),
    .B1(_3036_),
    .B2(_2996_),
    .ZN(_3037_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7788_ (.I(_0350_),
    .Z(_3038_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7789_ (.A1(_3009_),
    .A2(_2786_),
    .B(_3038_),
    .ZN(_3039_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7790_ (.A1(_2526_),
    .A2(_3037_),
    .B(_3039_),
    .ZN(_0182_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7791_ (.A1(\as2650.pc[11] ),
    .A2(_1657_),
    .Z(_3040_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7792_ (.A1(_2999_),
    .A2(_1142_),
    .ZN(_3041_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7793_ (.A1(_3015_),
    .A2(_3019_),
    .B(_3041_),
    .ZN(_3042_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7794_ (.A1(_3040_),
    .A2(_3042_),
    .ZN(_3043_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7795_ (.I(\as2650.addr_buff[3] ),
    .ZN(_3044_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7796_ (.I(_3044_),
    .Z(_3045_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7797_ (.A1(_3045_),
    .A2(_3003_),
    .Z(_3046_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7798_ (.A1(_3045_),
    .A2(_3006_),
    .Z(_3047_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7799_ (.A1(_2566_),
    .A2(_3046_),
    .B1(_3047_),
    .B2(_2744_),
    .ZN(_3048_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7800_ (.I(net40),
    .Z(_3049_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7801_ (.I(net39),
    .ZN(_3050_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7802_ (.A1(_3050_),
    .A2(_3010_),
    .ZN(_3051_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7803_ (.A1(_3049_),
    .A2(_3051_),
    .ZN(_3052_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7804_ (.A1(_2678_),
    .A2(_3048_),
    .B1(_3052_),
    .B2(_2620_),
    .C(_0417_),
    .ZN(_3053_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7805_ (.A1(_0418_),
    .A2(_3043_),
    .B(_3053_),
    .ZN(_3054_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7806_ (.A1(_3015_),
    .A2(_3023_),
    .B(_3041_),
    .ZN(_3055_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7807_ (.A1(_3040_),
    .A2(_3055_),
    .Z(_3056_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7808_ (.A1(_2537_),
    .A2(_3056_),
    .ZN(_3057_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7809_ (.A1(_3049_),
    .A2(_2542_),
    .B(_3057_),
    .ZN(_3058_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7810_ (.A1(_2550_),
    .A2(_3044_),
    .ZN(_3059_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7811_ (.A1(_3049_),
    .A2(_4431_),
    .B(_2721_),
    .C(_3059_),
    .ZN(_3060_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7812_ (.A1(_2553_),
    .A2(_3052_),
    .B(_3060_),
    .C(_2989_),
    .ZN(_3061_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7813_ (.A1(_1408_),
    .A2(_0377_),
    .B(_3061_),
    .ZN(_3062_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7814_ (.A1(_2886_),
    .A2(_3058_),
    .B1(_3062_),
    .B2(_4406_),
    .ZN(_3063_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7815_ (.A1(_1409_),
    .A2(_2959_),
    .B1(_3063_),
    .B2(_2993_),
    .ZN(_3064_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7816_ (.A1(_2814_),
    .A2(_3054_),
    .B1(_3064_),
    .B2(_2961_),
    .ZN(_3065_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7817_ (.A1(_1409_),
    .A2(_2530_),
    .B1(_3065_),
    .B2(_2996_),
    .ZN(_3066_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7818_ (.A1(_3049_),
    .A2(_2786_),
    .B(_3038_),
    .ZN(_3067_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7819_ (.A1(_2526_),
    .A2(_3066_),
    .B(_3067_),
    .ZN(_0183_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7820_ (.I(\as2650.pc[12] ),
    .Z(_3068_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7821_ (.I(_3068_),
    .Z(_3069_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7822_ (.I(\as2650.addr_buff[4] ),
    .Z(_3070_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7823_ (.A1(_3045_),
    .A2(_3006_),
    .ZN(_3071_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7824_ (.A1(_3070_),
    .A2(_3071_),
    .ZN(_3072_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7825_ (.A1(_3045_),
    .A2(_3003_),
    .ZN(_3073_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7826_ (.A1(_3070_),
    .A2(_3073_),
    .ZN(_3074_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7827_ (.A1(_2686_),
    .A2(_3072_),
    .B1(_3074_),
    .B2(_2929_),
    .ZN(_3075_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7828_ (.A1(net40),
    .A2(_3051_),
    .ZN(_3076_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7829_ (.A1(net53),
    .A2(_3076_),
    .Z(_3077_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7830_ (.A1(_2808_),
    .A2(_3077_),
    .ZN(_3078_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7831_ (.A1(_2795_),
    .A2(_3075_),
    .B(_3078_),
    .C(_2700_),
    .ZN(_3079_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7832_ (.A1(_3014_),
    .A2(_3040_),
    .ZN(_3080_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7833_ (.A1(_1406_),
    .A2(_1142_),
    .ZN(_3081_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7834_ (.A1(_3041_),
    .A2(_3016_),
    .A3(_3081_),
    .ZN(_3082_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7835_ (.A1(_3018_),
    .A2(_3080_),
    .B(_3082_),
    .ZN(_3083_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7836_ (.A1(\as2650.pc[12] ),
    .A2(_1142_),
    .Z(_3084_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7837_ (.A1(_3083_),
    .A2(_3084_),
    .ZN(_3085_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7838_ (.A1(_4410_),
    .A2(_3085_),
    .B(_2943_),
    .ZN(_3086_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7839_ (.A1(_3022_),
    .A2(_3080_),
    .B(_3082_),
    .ZN(_3087_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7840_ (.A1(_3084_),
    .A2(_3087_),
    .Z(_3088_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7841_ (.A1(_2537_),
    .A2(_3088_),
    .ZN(_3089_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7842_ (.A1(net53),
    .A2(_2542_),
    .B(_3089_),
    .ZN(_3090_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7843_ (.A1(_2768_),
    .A2(_3070_),
    .ZN(_3091_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7844_ (.A1(net53),
    .A2(_2821_),
    .B(_2721_),
    .ZN(_3092_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _7845_ (.A1(_4436_),
    .A2(_3077_),
    .B1(_3091_),
    .B2(_3092_),
    .C(_2989_),
    .ZN(_3093_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7846_ (.A1(_3069_),
    .A2(_2531_),
    .B(_3093_),
    .ZN(_3094_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7847_ (.A1(_2886_),
    .A2(_3090_),
    .B1(_3094_),
    .B2(_4406_),
    .ZN(_3095_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7848_ (.A1(_3069_),
    .A2(_2959_),
    .B1(_3095_),
    .B2(_2861_),
    .ZN(_3096_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7849_ (.A1(_3079_),
    .A2(_3086_),
    .B1(_3096_),
    .B2(_0306_),
    .ZN(_3097_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7850_ (.A1(_3069_),
    .A2(_2530_),
    .B1(_3097_),
    .B2(_2996_),
    .ZN(_3098_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7851_ (.A1(net53),
    .A2(_2786_),
    .B(_3038_),
    .ZN(_3099_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7852_ (.A1(_2526_),
    .A2(_3098_),
    .B(_3099_),
    .ZN(_0184_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7853_ (.A1(_4222_),
    .A2(_1482_),
    .A3(_0557_),
    .ZN(_3100_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _7854_ (.A1(_2511_),
    .A2(_2517_),
    .Z(_3101_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7855_ (.A1(_1626_),
    .A2(_1247_),
    .ZN(_3102_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7856_ (.A1(_4334_),
    .A2(_2492_),
    .A3(_2494_),
    .ZN(_3103_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _7857_ (.A1(_4337_),
    .A2(_0330_),
    .A3(_3103_),
    .ZN(_3104_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _7858_ (.A1(_2555_),
    .A2(_0420_),
    .A3(_1482_),
    .A4(_2344_),
    .Z(_3105_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _7859_ (.A1(_2487_),
    .A2(_3102_),
    .A3(_3104_),
    .A4(_3105_),
    .ZN(_3106_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _7860_ (.A1(_0423_),
    .A2(_4402_),
    .A3(_4256_),
    .A4(_2486_),
    .ZN(_3107_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7861_ (.A1(_2489_),
    .A2(_2499_),
    .ZN(_3108_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7862_ (.I(_2512_),
    .ZN(_3109_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7863_ (.A1(_4416_),
    .A2(_0315_),
    .B(_2495_),
    .ZN(_3110_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7864_ (.A1(_1481_),
    .A2(_0552_),
    .ZN(_3111_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _7865_ (.A1(_0411_),
    .A2(_2712_),
    .A3(_3111_),
    .ZN(_3112_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _7866_ (.A1(_3109_),
    .A2(_2496_),
    .A3(_3110_),
    .A4(_3112_),
    .ZN(_3113_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _7867_ (.A1(_3106_),
    .A2(_3107_),
    .A3(_3108_),
    .A4(_3113_),
    .ZN(_3114_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7868_ (.A1(_3101_),
    .A2(_3114_),
    .ZN(_3115_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7869_ (.A1(_2507_),
    .A2(_3100_),
    .A3(_3115_),
    .ZN(_3116_));
 gf180mcu_fd_sc_mcu7t5v0__oai222_1 _7870_ (.A1(_0386_),
    .A2(_0442_),
    .B1(_0361_),
    .B2(_0454_),
    .C1(_0303_),
    .C2(net27),
    .ZN(_3117_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7871_ (.A1(_2673_),
    .A2(_1525_),
    .B1(_3117_),
    .B2(_1252_),
    .ZN(_3118_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7872_ (.A1(_3116_),
    .A2(_3118_),
    .ZN(_3119_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7873_ (.A1(net50),
    .A2(_3116_),
    .B(_3119_),
    .C(_2629_),
    .ZN(_0185_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7874_ (.A1(_0434_),
    .A2(_2518_),
    .ZN(_3120_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _7875_ (.A1(_4267_),
    .A2(_4275_),
    .A3(_2518_),
    .ZN(_3121_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _7876_ (.A1(_3120_),
    .A2(_3102_),
    .A3(_3121_),
    .ZN(_3122_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _7877_ (.A1(_0342_),
    .A2(_4241_),
    .A3(_1252_),
    .ZN(_3123_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _7878_ (.A1(_4405_),
    .A2(_0345_),
    .A3(_2518_),
    .ZN(_3124_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7879_ (.A1(_0311_),
    .A2(_3123_),
    .B(_3124_),
    .ZN(_3125_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7880_ (.A1(_4048_),
    .A2(_4415_),
    .ZN(_3126_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _7881_ (.A1(_2498_),
    .A2(_3126_),
    .A3(_2342_),
    .ZN(_3127_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7882_ (.I(_2352_),
    .Z(_3128_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7883_ (.A1(_0310_),
    .A2(_2494_),
    .ZN(_3129_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7884_ (.A1(_3128_),
    .A2(_3111_),
    .B(_3129_),
    .ZN(_3130_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _7885_ (.A1(_0432_),
    .A2(_2487_),
    .A3(_3127_),
    .A4(_3130_),
    .ZN(_3131_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7886_ (.I(_0360_),
    .Z(_3132_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _7887_ (.A1(_1258_),
    .A2(_0430_),
    .A3(_0679_),
    .ZN(_3133_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _7888_ (.A1(_0385_),
    .A2(_3132_),
    .A3(_2486_),
    .A4(_3133_),
    .ZN(_3134_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7889_ (.A1(_3108_),
    .A2(_3131_),
    .A3(_3134_),
    .ZN(_3135_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7890_ (.A1(_3101_),
    .A2(_3135_),
    .ZN(_3136_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _7891_ (.A1(_2503_),
    .A2(_3122_),
    .A3(_3125_),
    .A4(_3136_),
    .ZN(_3137_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7892_ (.A1(_2500_),
    .A2(_3137_),
    .ZN(_3138_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7893_ (.I(_4423_),
    .Z(_3139_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7894_ (.A1(_4262_),
    .A2(_2334_),
    .ZN(_3140_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7895_ (.A1(_3139_),
    .A2(_4428_),
    .B(_2600_),
    .C(_4432_),
    .ZN(_3141_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _7896_ (.A1(_3139_),
    .A2(_4349_),
    .A3(_3140_),
    .B(_3141_),
    .ZN(_3142_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7897_ (.A1(net52),
    .A2(_3142_),
    .B(_0414_),
    .ZN(_3143_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7898_ (.A1(_2385_),
    .A2(_0415_),
    .B(_3143_),
    .C(_0438_),
    .ZN(_3144_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7899_ (.A1(net52),
    .A2(_0299_),
    .A3(_0380_),
    .ZN(_3145_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7900_ (.A1(net52),
    .A2(_0321_),
    .A3(_1519_),
    .ZN(_3146_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _7901_ (.A1(_0381_),
    .A2(_3145_),
    .B1(_3146_),
    .B2(_4349_),
    .C(_2486_),
    .ZN(_3147_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7902_ (.A1(_0309_),
    .A2(_1749_),
    .ZN(_3148_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7903_ (.A1(_3144_),
    .A2(_3147_),
    .B(_3148_),
    .ZN(_3149_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7904_ (.A1(net52),
    .A2(_3138_),
    .ZN(_3150_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7905_ (.A1(_3138_),
    .A2(_3149_),
    .B(_3150_),
    .C(_2629_),
    .ZN(_0186_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7906_ (.A1(_0313_),
    .A2(_0327_),
    .ZN(_3151_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7907_ (.A1(_0299_),
    .A2(_2492_),
    .A3(_3151_),
    .ZN(_3152_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7908_ (.A1(_1588_),
    .A2(_3152_),
    .ZN(_3153_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7909_ (.A1(_0315_),
    .A2(_2495_),
    .ZN(_3154_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _7910_ (.A1(_2504_),
    .A2(_2512_),
    .A3(_2513_),
    .ZN(_3155_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _7911_ (.A1(_1482_),
    .A2(_3153_),
    .B(_3154_),
    .C(_3155_),
    .ZN(_3156_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7912_ (.A1(_2380_),
    .A2(_2478_),
    .ZN(_3157_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7913_ (.A1(_0597_),
    .A2(_3156_),
    .ZN(_3158_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7914_ (.A1(_3156_),
    .A2(_3157_),
    .B(_3158_),
    .C(_2629_),
    .ZN(_0187_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7915_ (.A1(_2382_),
    .A2(_2478_),
    .ZN(_3159_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7916_ (.A1(_0596_),
    .A2(_3156_),
    .ZN(_3160_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7917_ (.I(_1507_),
    .Z(_3161_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7918_ (.A1(_3156_),
    .A2(_3159_),
    .B(_3160_),
    .C(_3161_),
    .ZN(_0188_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7919_ (.I(_1259_),
    .Z(_3162_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7920_ (.A1(_0490_),
    .A2(_0497_),
    .B(_0369_),
    .ZN(_3163_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7921_ (.A1(_1463_),
    .A2(_3163_),
    .ZN(_3164_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _7922_ (.A1(_1802_),
    .A2(_3162_),
    .A3(_0530_),
    .A4(_3164_),
    .ZN(_3165_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7923_ (.I(_3165_),
    .Z(_3166_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7924_ (.A1(_0663_),
    .A2(_1463_),
    .ZN(_3167_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7925_ (.I(_4047_),
    .Z(_3168_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7926_ (.I(_3168_),
    .Z(_3169_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7927_ (.I(_3169_),
    .Z(_3170_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7928_ (.A1(_3170_),
    .A2(_1676_),
    .ZN(_3171_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7929_ (.A1(_3167_),
    .A2(_3171_),
    .ZN(_3172_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7930_ (.A1(_3166_),
    .A2(_3172_),
    .ZN(_3173_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7931_ (.A1(_0584_),
    .A2(_3166_),
    .B(_3173_),
    .ZN(_0189_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7932_ (.I(_2473_),
    .Z(_3174_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7933_ (.I(_2407_),
    .Z(_3175_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7934_ (.I(_3175_),
    .Z(_3176_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7935_ (.A1(_1540_),
    .A2(_3176_),
    .ZN(_3177_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7936_ (.A1(_3174_),
    .A2(_2365_),
    .B(_3177_),
    .ZN(_3178_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7937_ (.I0(_3178_),
    .I1(\as2650.holding_reg[1] ),
    .S(_3166_),
    .Z(_3179_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7938_ (.I(_3179_),
    .Z(_0190_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7939_ (.A1(_1545_),
    .A2(_1499_),
    .ZN(_3180_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7940_ (.A1(_3170_),
    .A2(_1678_),
    .ZN(_3181_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7941_ (.A1(_3180_),
    .A2(_3181_),
    .ZN(_3182_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7942_ (.I0(_3182_),
    .I1(\as2650.holding_reg[2] ),
    .S(_3166_),
    .Z(_3183_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7943_ (.I(_3183_),
    .Z(_0191_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7944_ (.A1(_4362_),
    .A2(_1680_),
    .ZN(_3184_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _7945_ (.A1(_0970_),
    .A2(_3174_),
    .B(_3184_),
    .ZN(_3185_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7946_ (.I(_3165_),
    .Z(_3186_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7947_ (.I0(_3185_),
    .I1(\as2650.holding_reg[3] ),
    .S(_3186_),
    .Z(_3187_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7948_ (.I(_3187_),
    .Z(_0192_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7949_ (.I(_3170_),
    .Z(_3188_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7950_ (.A1(_3188_),
    .A2(_2377_),
    .ZN(_3189_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7951_ (.A1(_1018_),
    .A2(_3176_),
    .ZN(_3190_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7952_ (.A1(_3189_),
    .A2(_3190_),
    .ZN(_3191_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7953_ (.I0(_3191_),
    .I1(\as2650.holding_reg[4] ),
    .S(_3186_),
    .Z(_3192_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7954_ (.I(_3192_),
    .Z(_0193_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7955_ (.I0(_1503_),
    .I1(_1056_),
    .S(_3186_),
    .Z(_3193_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7956_ (.I(_3193_),
    .Z(_0194_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7957_ (.I(_2407_),
    .Z(_3194_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7958_ (.I(_3194_),
    .Z(_3195_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7959_ (.A1(_3195_),
    .A2(_1674_),
    .ZN(_3196_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7960_ (.A1(_1122_),
    .A2(_3174_),
    .B(_3196_),
    .ZN(_3197_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7961_ (.I0(_3197_),
    .I1(\as2650.holding_reg[6] ),
    .S(_3186_),
    .Z(_3198_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7962_ (.I(_3198_),
    .Z(_0195_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7963_ (.A1(_1737_),
    .A2(_3126_),
    .ZN(_3199_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7964_ (.I0(_3199_),
    .I1(\as2650.holding_reg[7] ),
    .S(_3165_),
    .Z(_3200_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7965_ (.I(_3200_),
    .Z(_0196_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7966_ (.A1(_4450_),
    .A2(_4399_),
    .A3(_1279_),
    .ZN(_3201_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7967_ (.I(_0469_),
    .Z(_3202_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7968_ (.A1(_0336_),
    .A2(_3201_),
    .B(_3202_),
    .ZN(_0197_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7969_ (.I(\as2650.psu[7] ),
    .ZN(_3203_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7970_ (.A1(_0472_),
    .A2(_1694_),
    .B(_1495_),
    .C(_1654_),
    .ZN(_3204_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7971_ (.A1(_3203_),
    .A2(_0394_),
    .B(_3204_),
    .ZN(_3205_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7972_ (.A1(_3111_),
    .A2(_3205_),
    .B(net4),
    .C(_2510_),
    .ZN(_3206_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7973_ (.I(_2510_),
    .ZN(_3207_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7974_ (.A1(_1655_),
    .A2(_1722_),
    .ZN(_3208_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _7975_ (.A1(_0300_),
    .A2(_2498_),
    .A3(_3208_),
    .ZN(_3209_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7976_ (.A1(_1240_),
    .A2(_3207_),
    .B1(_3205_),
    .B2(_3209_),
    .C(_0465_),
    .ZN(_3210_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7977_ (.A1(_3203_),
    .A2(_0433_),
    .B1(_3206_),
    .B2(_3210_),
    .C(_0334_),
    .ZN(_0198_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7978_ (.A1(_0403_),
    .A2(_2495_),
    .B(_3103_),
    .C(_2480_),
    .ZN(_3211_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7979_ (.I(_3211_),
    .ZN(_3212_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _7980_ (.A1(_4384_),
    .A2(_1266_),
    .B1(_2488_),
    .B2(_4327_),
    .C(_3212_),
    .ZN(_3213_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7981_ (.A1(_2497_),
    .A2(_2501_),
    .ZN(_3214_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7982_ (.A1(_3122_),
    .A2(_3125_),
    .ZN(_3215_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _7983_ (.A1(_3155_),
    .A2(_3213_),
    .A3(_3214_),
    .A4(_3215_),
    .ZN(_3216_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _7984_ (.A1(_2768_),
    .A2(_4241_),
    .A3(_2863_),
    .B(_4286_),
    .ZN(_3217_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7985_ (.A1(_2519_),
    .A2(_3217_),
    .B(_3101_),
    .ZN(_3218_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7986_ (.A1(_3216_),
    .A2(_3218_),
    .ZN(_3219_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7987_ (.I(_3219_),
    .Z(_3220_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7988_ (.I(_2781_),
    .Z(_3221_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7989_ (.I(_1276_),
    .Z(_3222_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7990_ (.A1(_1275_),
    .A2(_0429_),
    .Z(_3223_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _7991_ (.A1(_1217_),
    .A2(_4188_),
    .A3(_4220_),
    .ZN(_3224_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7992_ (.I0(_3222_),
    .I1(_3223_),
    .S(_3224_),
    .Z(_3225_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7993_ (.I0(_3223_),
    .I1(_3222_),
    .S(_4236_),
    .Z(_3226_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7994_ (.I0(_3225_),
    .I1(_3226_),
    .S(_4057_),
    .Z(_3227_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7995_ (.A1(_1276_),
    .A2(_0392_),
    .ZN(_3228_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7996_ (.A1(_2715_),
    .A2(_2539_),
    .B(_3228_),
    .C(_0399_),
    .ZN(_3229_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7997_ (.A1(_3222_),
    .A2(_2596_),
    .B1(_0463_),
    .B2(_2329_),
    .C(_0814_),
    .ZN(_3230_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7998_ (.A1(_2362_),
    .A2(_3140_),
    .B(_3229_),
    .C(_3230_),
    .ZN(_3231_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7999_ (.I(_3132_),
    .Z(_3232_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8000_ (.A1(_4050_),
    .A2(_3227_),
    .B(_3231_),
    .C(_3232_),
    .ZN(_3233_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8001_ (.A1(_2352_),
    .A2(_1259_),
    .ZN(_3234_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8002_ (.I(_3234_),
    .Z(_3235_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8003_ (.A1(_4161_),
    .A2(_2891_),
    .ZN(_3236_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8004_ (.A1(_1676_),
    .A2(_3236_),
    .Z(_3237_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8005_ (.I(_3128_),
    .Z(_3238_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8006_ (.A1(_3238_),
    .A2(_2331_),
    .ZN(_3239_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8007_ (.A1(_3235_),
    .A2(_3237_),
    .B1(_3239_),
    .B2(_1277_),
    .C(_3033_),
    .ZN(_3240_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8008_ (.I(_2454_),
    .Z(_3241_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8009_ (.I(_3241_),
    .Z(_3242_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8010_ (.A1(_0699_),
    .A2(_0701_),
    .ZN(_3243_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8011_ (.I(_3243_),
    .Z(_3244_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8012_ (.I(_3244_),
    .Z(_3245_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8013_ (.I(_2387_),
    .Z(_3246_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _8014_ (.A1(\as2650.stack[3][0] ),
    .A2(_3246_),
    .B1(_1573_),
    .B2(\as2650.stack[2][0] ),
    .ZN(_3247_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _8015_ (.I(_3247_),
    .ZN(_3248_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _8016_ (.A1(\as2650.stack[1][0] ),
    .A2(_3242_),
    .B1(_3245_),
    .B2(\as2650.stack[0][0] ),
    .C(_3248_),
    .ZN(_3249_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8017_ (.I(_2387_),
    .Z(_3250_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8018_ (.I(_1572_),
    .Z(_3251_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8019_ (.I(_3241_),
    .Z(_3252_));
 gf180mcu_fd_sc_mcu7t5v0__oai222_1 _8020_ (.A1(\as2650.stack[7][0] ),
    .A2(_3250_),
    .B1(_3251_),
    .B2(\as2650.stack[6][0] ),
    .C1(_3252_),
    .C2(\as2650.stack[5][0] ),
    .ZN(_3253_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8021_ (.I(_3244_),
    .Z(_3254_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8022_ (.A1(\as2650.stack[4][0] ),
    .A2(_3254_),
    .B(_0906_),
    .ZN(_3255_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _8023_ (.A1(_0973_),
    .A2(_3249_),
    .B1(_3253_),
    .B2(_3255_),
    .ZN(_3256_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8024_ (.I(_4301_),
    .Z(_3257_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8025_ (.I(_3257_),
    .Z(_3258_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8026_ (.A1(_1693_),
    .A2(_2539_),
    .B(_3228_),
    .C(_3169_),
    .ZN(_3259_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8027_ (.I(_2471_),
    .Z(_3260_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8028_ (.A1(_3222_),
    .A2(_3260_),
    .ZN(_3261_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8029_ (.A1(_0414_),
    .A2(_3259_),
    .A3(_3261_),
    .ZN(_3262_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8030_ (.A1(_1509_),
    .A2(_0338_),
    .ZN(_3263_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8031_ (.A1(_1277_),
    .A2(_1511_),
    .B(_3262_),
    .C(_3263_),
    .ZN(_3264_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8032_ (.A1(_3233_),
    .A2(_3240_),
    .B1(_3256_),
    .B2(_3258_),
    .C(_3264_),
    .ZN(_3265_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8033_ (.A1(_2527_),
    .A2(_3221_),
    .B(_3265_),
    .ZN(_3266_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8034_ (.A1(_3220_),
    .A2(_3266_),
    .ZN(_3267_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _8035_ (.A1(_3216_),
    .A2(_3218_),
    .Z(_3268_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8036_ (.I(_3268_),
    .Z(_3269_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8037_ (.A1(_2527_),
    .A2(_3269_),
    .B(_1687_),
    .ZN(_3270_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8038_ (.A1(_3267_),
    .A2(_3270_),
    .ZN(_0199_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8039_ (.I(_3219_),
    .Z(_3271_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8040_ (.I(_3271_),
    .Z(_3272_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8041_ (.I(_3263_),
    .Z(_3273_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8042_ (.A1(_1287_),
    .A2(_1275_),
    .Z(_3274_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8043_ (.I(_3274_),
    .Z(_3275_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8044_ (.A1(_4221_),
    .A2(_4237_),
    .B(_0812_),
    .ZN(_3276_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8045_ (.A1(_4423_),
    .A2(_3276_),
    .ZN(_3277_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8046_ (.I(_3277_),
    .Z(_3278_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8047_ (.A1(_1274_),
    .A2(_4268_),
    .ZN(_3279_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8048_ (.A1(_2582_),
    .A2(_3279_),
    .Z(_3280_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _8049_ (.A1(_3168_),
    .A2(_4222_),
    .A3(_4237_),
    .B1(_0388_),
    .B2(_2330_),
    .ZN(_3281_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8050_ (.I(_3281_),
    .Z(_3282_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _8051_ (.A1(net7),
    .A2(_4161_),
    .Z(_3283_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8052_ (.A1(_0784_),
    .A2(_4151_),
    .Z(_3284_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8053_ (.A1(_3283_),
    .A2(_3284_),
    .B(_4448_),
    .ZN(_3285_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8054_ (.A1(_3283_),
    .A2(_3284_),
    .B(_3285_),
    .ZN(_3286_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8055_ (.A1(_0787_),
    .A2(_2334_),
    .ZN(_3287_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8056_ (.A1(_2353_),
    .A2(_3286_),
    .A3(_3287_),
    .ZN(_3288_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8057_ (.A1(_2263_),
    .A2(_2590_),
    .ZN(_3289_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8058_ (.A1(_1287_),
    .A2(_2536_),
    .B(_3289_),
    .ZN(_3290_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8059_ (.A1(_0398_),
    .A2(_3290_),
    .ZN(_3291_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8060_ (.I(_0462_),
    .Z(_3292_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8061_ (.A1(_4345_),
    .A2(_4434_),
    .ZN(_3293_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8062_ (.A1(_0375_),
    .A2(_3274_),
    .ZN(_3294_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8063_ (.A1(_0787_),
    .A2(_3292_),
    .B1(_3293_),
    .B2(_2366_),
    .C(_3294_),
    .ZN(_3295_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8064_ (.A1(_0360_),
    .A2(_3291_),
    .A3(_3295_),
    .ZN(_3296_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8065_ (.A1(_3288_),
    .A2(_3296_),
    .B(_0814_),
    .ZN(_3297_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _8066_ (.A1(_3032_),
    .A2(_3297_),
    .Z(_3298_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8067_ (.A1(_3278_),
    .A2(_3280_),
    .B1(_3275_),
    .B2(_3282_),
    .C(_3298_),
    .ZN(_3299_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8068_ (.A1(_3175_),
    .A2(_3290_),
    .B(_0414_),
    .ZN(_3300_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8069_ (.A1(_4362_),
    .A2(_3275_),
    .B(_3300_),
    .ZN(_3301_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8070_ (.I(_3246_),
    .Z(_3302_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8071_ (.I(_1573_),
    .Z(_3303_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _8072_ (.A1(\as2650.stack[7][1] ),
    .A2(_3302_),
    .B1(_3303_),
    .B2(\as2650.stack[6][1] ),
    .ZN(_3304_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _8073_ (.A1(\as2650.stack[5][1] ),
    .A2(_2456_),
    .B1(_3254_),
    .B2(\as2650.stack[4][1] ),
    .C(_0906_),
    .ZN(_3305_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _8074_ (.A1(\as2650.stack[3][1] ),
    .A2(_3302_),
    .B1(_3303_),
    .B2(\as2650.stack[2][1] ),
    .ZN(_3306_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _8075_ (.A1(\as2650.stack[1][1] ),
    .A2(_3242_),
    .B1(_3254_),
    .B2(\as2650.stack[0][1] ),
    .C(_0722_),
    .ZN(_3307_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _8076_ (.A1(_3304_),
    .A2(_3305_),
    .B1(_3306_),
    .B2(_3307_),
    .ZN(_3308_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8077_ (.A1(_1510_),
    .A2(_3308_),
    .ZN(_3309_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8078_ (.I(_4367_),
    .Z(_3310_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8079_ (.A1(_1510_),
    .A2(_3275_),
    .B(_3309_),
    .C(_3310_),
    .ZN(_3311_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _8080_ (.A1(_3299_),
    .A2(_3301_),
    .A3(_3311_),
    .B(_3273_),
    .ZN(_3312_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8081_ (.I(_3268_),
    .Z(_3313_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8082_ (.A1(_3273_),
    .A2(_3275_),
    .B(_3312_),
    .C(_3313_),
    .ZN(_3314_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8083_ (.A1(_1687_),
    .A2(_3314_),
    .ZN(_3315_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8084_ (.A1(_1288_),
    .A2(_3272_),
    .B(_3315_),
    .ZN(_0200_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8085_ (.I(_2731_),
    .Z(_3316_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8086_ (.A1(_2582_),
    .A2(_1275_),
    .ZN(_3317_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _8087_ (.A1(_2664_),
    .A2(_3317_),
    .ZN(_3318_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8088_ (.A1(_1716_),
    .A2(_4135_),
    .Z(_3319_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _8089_ (.A1(_0785_),
    .A2(_4151_),
    .Z(_3320_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8090_ (.A1(_3283_),
    .A2(_3284_),
    .B(_3320_),
    .ZN(_3321_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8091_ (.A1(_3319_),
    .A2(_3321_),
    .Z(_3322_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8092_ (.A1(_3027_),
    .A2(_3322_),
    .ZN(_3323_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8093_ (.A1(_2369_),
    .A2(_2666_),
    .B(_3323_),
    .ZN(_3324_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8094_ (.A1(_2663_),
    .A2(_1692_),
    .ZN(_3325_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8095_ (.A1(_2586_),
    .A2(_2660_),
    .B(_3325_),
    .ZN(_3326_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8096_ (.A1(_2663_),
    .A2(_3317_),
    .Z(_3327_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8097_ (.A1(\as2650.addr_buff[2] ),
    .A2(_3140_),
    .ZN(_3328_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8098_ (.A1(_2369_),
    .A2(_3292_),
    .B1(_3327_),
    .B2(_2596_),
    .C(_3328_),
    .ZN(_3329_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8099_ (.A1(_2713_),
    .A2(_3326_),
    .B(_3329_),
    .ZN(_3330_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8100_ (.A1(_3132_),
    .A2(_3330_),
    .ZN(_3331_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8101_ (.A1(_4429_),
    .A2(_3324_),
    .B(_3331_),
    .ZN(_3332_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8102_ (.A1(_4050_),
    .A2(_3332_),
    .ZN(_3333_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8103_ (.A1(_0436_),
    .A2(_3333_),
    .ZN(_3334_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8104_ (.A1(_1287_),
    .A2(_3279_),
    .ZN(_3335_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _8105_ (.A1(_2664_),
    .A2(_3335_),
    .ZN(_3336_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8106_ (.A1(_3278_),
    .A2(_3336_),
    .B1(_3327_),
    .B2(_3282_),
    .ZN(_3337_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _8107_ (.I(_3337_),
    .ZN(_3338_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8108_ (.I(_1474_),
    .Z(_3339_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8109_ (.A1(_1489_),
    .A2(_3327_),
    .ZN(_3340_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8110_ (.A1(_3339_),
    .A2(_3326_),
    .B(_3340_),
    .C(_0415_),
    .ZN(_3341_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8111_ (.A1(_3334_),
    .A2(_3338_),
    .B(_3341_),
    .C(_0424_),
    .ZN(_3342_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8112_ (.A1(_4294_),
    .A2(_0445_),
    .ZN(_3343_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8113_ (.I(_3343_),
    .Z(_3344_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _8114_ (.A1(\as2650.stack[7][2] ),
    .A2(_3250_),
    .B1(_3251_),
    .B2(\as2650.stack[6][2] ),
    .ZN(_3345_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _8115_ (.A1(\as2650.stack[5][2] ),
    .A2(_3252_),
    .B1(_3245_),
    .B2(\as2650.stack[4][2] ),
    .C(_0905_),
    .ZN(_3346_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8116_ (.I(_1572_),
    .Z(_3347_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _8117_ (.A1(\as2650.stack[3][2] ),
    .A2(_2388_),
    .B1(_3347_),
    .B2(\as2650.stack[2][2] ),
    .ZN(_3348_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _8118_ (.A1(\as2650.stack[1][2] ),
    .A2(_3252_),
    .B1(_3245_),
    .B2(\as2650.stack[0][2] ),
    .C(_1046_),
    .ZN(_3349_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _8119_ (.A1(_3345_),
    .A2(_3346_),
    .B1(_3348_),
    .B2(_3349_),
    .ZN(_3350_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _8120_ (.I(_3350_),
    .ZN(_3351_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8121_ (.A1(_3344_),
    .A2(_3327_),
    .B1(_3351_),
    .B2(_3258_),
    .C(_2816_),
    .ZN(_3352_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8122_ (.A1(_3316_),
    .A2(_3318_),
    .B1(_3342_),
    .B2(_3352_),
    .C(_3220_),
    .ZN(_3353_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8123_ (.I(_1686_),
    .Z(_3354_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8124_ (.A1(_2664_),
    .A2(_3269_),
    .B(_3354_),
    .ZN(_3355_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8125_ (.A1(_3353_),
    .A2(_3355_),
    .ZN(_0201_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _8126_ (.A1(\as2650.pc[2] ),
    .A2(_2582_),
    .A3(_1274_),
    .ZN(_3356_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8127_ (.A1(_1298_),
    .A2(_3356_),
    .Z(_3357_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _8128_ (.I(_3282_),
    .ZN(_3358_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _8129_ (.A1(_2663_),
    .A2(_3335_),
    .ZN(_3359_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8130_ (.A1(_2710_),
    .A2(_3359_),
    .Z(_3360_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _8131_ (.A1(_0952_),
    .A2(_4130_),
    .Z(_3361_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8132_ (.A1(_0952_),
    .A2(_4130_),
    .ZN(_3362_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _8133_ (.A1(_3361_),
    .A2(_3362_),
    .Z(_3363_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8134_ (.A1(_0881_),
    .A2(_4135_),
    .ZN(_3364_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8135_ (.A1(_3319_),
    .A2(_3321_),
    .B(_3364_),
    .ZN(_3365_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8136_ (.A1(_3363_),
    .A2(_3365_),
    .Z(_3366_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8137_ (.A1(_1680_),
    .A2(_2863_),
    .ZN(_3367_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8138_ (.A1(_2864_),
    .A2(_3366_),
    .B(_3367_),
    .C(_2354_),
    .ZN(_3368_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8139_ (.A1(_2710_),
    .A2(_3356_),
    .Z(_3369_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8140_ (.I(_3293_),
    .Z(_3370_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8141_ (.A1(_2263_),
    .A2(_2717_),
    .ZN(_3371_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8142_ (.A1(_1297_),
    .A2(_1216_),
    .B(_3371_),
    .ZN(_3372_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _8143_ (.A1(_1679_),
    .A2(_3292_),
    .B1(_3370_),
    .B2(\as2650.addr_buff[3] ),
    .C1(_3372_),
    .C2(_0398_),
    .ZN(_3373_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8144_ (.A1(_0376_),
    .A2(_3369_),
    .B(_3373_),
    .C(_3128_),
    .ZN(_3374_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8145_ (.A1(_3368_),
    .A2(_3374_),
    .B(_3260_),
    .ZN(_3375_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8146_ (.A1(_3277_),
    .A2(_3360_),
    .B(_3375_),
    .C(_3032_),
    .ZN(_3376_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8147_ (.A1(_3358_),
    .A2(_3357_),
    .B(_3376_),
    .ZN(_3377_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8148_ (.I(_3343_),
    .Z(_3378_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8149_ (.I(_3243_),
    .Z(_3379_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8150_ (.I(_3379_),
    .Z(_3380_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _8151_ (.A1(\as2650.stack[5][3] ),
    .A2(_2455_),
    .B1(_3347_),
    .B2(\as2650.stack[6][3] ),
    .ZN(_3381_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _8152_ (.I(_3381_),
    .ZN(_3382_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _8153_ (.A1(\as2650.stack[7][3] ),
    .A2(_2389_),
    .B1(_3380_),
    .B2(\as2650.stack[4][3] ),
    .C(_3382_),
    .ZN(_3383_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _8154_ (.A1(\as2650.stack[3][3] ),
    .A2(_3302_),
    .B1(_1574_),
    .B2(\as2650.stack[2][3] ),
    .ZN(_3384_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _8155_ (.A1(\as2650.stack[1][3] ),
    .A2(_2456_),
    .B1(_3254_),
    .B2(\as2650.stack[0][3] ),
    .C(_0825_),
    .ZN(_3385_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _8156_ (.A1(_0831_),
    .A2(_3383_),
    .B1(_3384_),
    .B2(_3385_),
    .ZN(_3386_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8157_ (.A1(_2472_),
    .A2(_3372_),
    .ZN(_3387_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8158_ (.A1(_1474_),
    .A2(_3369_),
    .B(_3387_),
    .C(_0435_),
    .ZN(_3388_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8159_ (.A1(_3378_),
    .A2(_3357_),
    .B1(_3386_),
    .B2(_3257_),
    .C(_3388_),
    .ZN(_3389_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8160_ (.A1(_3377_),
    .A2(_3389_),
    .B(_2731_),
    .ZN(_3390_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8161_ (.I(_3219_),
    .Z(_3391_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8162_ (.A1(_3221_),
    .A2(_3357_),
    .B(_3390_),
    .C(_3391_),
    .ZN(_3392_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8163_ (.A1(_1298_),
    .A2(_3272_),
    .B(_3392_),
    .C(_3161_),
    .ZN(_0202_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8164_ (.A1(_1297_),
    .A2(_3356_),
    .ZN(_3393_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8165_ (.A1(_2767_),
    .A2(_3393_),
    .Z(_3394_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8166_ (.I(_3394_),
    .Z(_3395_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8167_ (.A1(_1297_),
    .A2(_3359_),
    .ZN(_3396_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8168_ (.A1(_1305_),
    .A2(_3396_),
    .Z(_3397_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _8169_ (.I(_3362_),
    .ZN(_3398_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8170_ (.A1(_3398_),
    .A2(_3365_),
    .B(_3361_),
    .ZN(_3399_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _8171_ (.A1(_1022_),
    .A2(_4120_),
    .A3(_3399_),
    .Z(_3400_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8172_ (.A1(_1672_),
    .A2(_2335_),
    .ZN(_3401_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8173_ (.A1(_2864_),
    .A2(_3400_),
    .B(_3401_),
    .C(_2354_),
    .ZN(_3402_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8174_ (.A1(_2596_),
    .A2(_3394_),
    .ZN(_3403_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8175_ (.A1(_2767_),
    .A2(_2585_),
    .ZN(_3404_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8176_ (.A1(_0391_),
    .A2(_2776_),
    .B(_3404_),
    .ZN(_3405_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _8177_ (.A1(_1023_),
    .A2(_3292_),
    .B1(_3370_),
    .B2(_3070_),
    .C1(_3405_),
    .C2(_0398_),
    .ZN(_3406_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8178_ (.A1(_3128_),
    .A2(_3403_),
    .A3(_3406_),
    .ZN(_3407_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8179_ (.A1(_3402_),
    .A2(_3407_),
    .ZN(_3408_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8180_ (.A1(_3277_),
    .A2(_3397_),
    .B1(_3408_),
    .B2(_3170_),
    .C(_3032_),
    .ZN(_3409_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8181_ (.A1(_3358_),
    .A2(_3395_),
    .B(_3409_),
    .ZN(_3410_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _8182_ (.A1(\as2650.stack[3][4] ),
    .A2(_2388_),
    .B1(_3347_),
    .B2(\as2650.stack[2][4] ),
    .ZN(_3411_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _8183_ (.A1(\as2650.stack[1][4] ),
    .A2(_3252_),
    .B1(_3379_),
    .B2(\as2650.stack[0][4] ),
    .C(_1046_),
    .ZN(_3412_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _8184_ (.A1(\as2650.stack[7][4] ),
    .A2(_2388_),
    .B1(_3347_),
    .B2(\as2650.stack[6][4] ),
    .ZN(_3413_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _8185_ (.A1(\as2650.stack[5][4] ),
    .A2(_2455_),
    .B1(_3379_),
    .B2(\as2650.stack[4][4] ),
    .C(_0905_),
    .ZN(_3414_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _8186_ (.A1(_3411_),
    .A2(_3412_),
    .B1(_3413_),
    .B2(_3414_),
    .ZN(_3415_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8187_ (.A1(_4049_),
    .A2(_3395_),
    .ZN(_3416_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8188_ (.A1(_4361_),
    .A2(_3405_),
    .B(_2548_),
    .ZN(_3417_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8189_ (.A1(_3416_),
    .A2(_3417_),
    .ZN(_3418_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8190_ (.A1(_3378_),
    .A2(_3395_),
    .B1(_3415_),
    .B2(_3257_),
    .C(_3418_),
    .ZN(_3419_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8191_ (.A1(_3410_),
    .A2(_3419_),
    .B(_2731_),
    .ZN(_3420_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8192_ (.A1(_3221_),
    .A2(_3395_),
    .B(_3420_),
    .C(_3391_),
    .ZN(_3421_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8193_ (.A1(_1305_),
    .A2(_3272_),
    .B(_3421_),
    .C(_3161_),
    .ZN(_0203_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8194_ (.I(_2781_),
    .Z(_3422_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _8195_ (.A1(_1304_),
    .A2(_1296_),
    .A3(_3356_),
    .ZN(_3423_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8196_ (.A1(_2789_),
    .A2(_3423_),
    .Z(_3424_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8197_ (.I(_3424_),
    .Z(_3425_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8198_ (.I(_3343_),
    .Z(_3426_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _8199_ (.A1(\as2650.stack[3][5] ),
    .A2(_3246_),
    .B1(_1573_),
    .B2(\as2650.stack[2][5] ),
    .ZN(_3427_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _8200_ (.A1(\as2650.stack[1][5] ),
    .A2(_2455_),
    .B1(_3379_),
    .B2(\as2650.stack[0][5] ),
    .C(_0721_),
    .ZN(_3428_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _8201_ (.A1(\as2650.stack[5][5] ),
    .A2(_3241_),
    .B1(_1572_),
    .B2(\as2650.stack[6][5] ),
    .ZN(_3429_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _8202_ (.I(_3429_),
    .ZN(_3430_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _8203_ (.A1(\as2650.stack[7][5] ),
    .A2(_3246_),
    .B1(_3244_),
    .B2(\as2650.stack[4][5] ),
    .C(_3430_),
    .ZN(_3431_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _8204_ (.A1(_3427_),
    .A2(_3428_),
    .B1(_3431_),
    .B2(_1046_),
    .ZN(_3432_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8205_ (.I(_3257_),
    .Z(_3433_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8206_ (.A1(_1314_),
    .A2(_4415_),
    .ZN(_3434_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8207_ (.A1(_2586_),
    .A2(_2819_),
    .B(_3434_),
    .ZN(_3435_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8208_ (.A1(_0737_),
    .A2(_0376_),
    .ZN(_3436_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8209_ (.A1(_0533_),
    .A2(_2334_),
    .ZN(_3437_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8210_ (.A1(_1501_),
    .A2(_4448_),
    .B(_3437_),
    .ZN(_3438_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8211_ (.A1(_3424_),
    .A2(_3436_),
    .B1(_3438_),
    .B2(_2330_),
    .ZN(_3439_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _8212_ (.A1(_0437_),
    .A2(_0679_),
    .A3(_3435_),
    .B(_3439_),
    .ZN(_3440_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8213_ (.I(_3276_),
    .Z(_3441_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _8214_ (.A1(_1313_),
    .A2(_1304_),
    .A3(_1296_),
    .A4(_3359_),
    .ZN(_3442_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8215_ (.A1(_2767_),
    .A2(_3396_),
    .B(_2789_),
    .ZN(_3443_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _8216_ (.A1(_3441_),
    .A2(_3442_),
    .A3(_3443_),
    .ZN(_3444_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8217_ (.A1(_3440_),
    .A2(_3444_),
    .B(_3132_),
    .ZN(_3445_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8218_ (.A1(_1019_),
    .A2(_4120_),
    .ZN(_3446_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8219_ (.A1(_1019_),
    .A2(_4120_),
    .ZN(_3447_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8220_ (.A1(_3446_),
    .A2(_3399_),
    .B(_3447_),
    .ZN(_3448_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _8221_ (.A1(_1500_),
    .A2(_4111_),
    .A3(_3448_),
    .Z(_3449_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8222_ (.A1(_1095_),
    .A2(_2552_),
    .B(_3234_),
    .ZN(_3450_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8223_ (.A1(_2723_),
    .A2(_3449_),
    .B(_3450_),
    .ZN(_3451_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8224_ (.A1(_3281_),
    .A2(_3425_),
    .B(_3451_),
    .C(_2548_),
    .ZN(_3452_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8225_ (.A1(_2407_),
    .A2(_3435_),
    .ZN(_3453_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8226_ (.A1(_3260_),
    .A2(_3425_),
    .B(_3453_),
    .ZN(_3454_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8227_ (.I(_4405_),
    .Z(_3455_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8228_ (.A1(_3445_),
    .A2(_3452_),
    .B1(_3454_),
    .B2(_3455_),
    .C(_2861_),
    .ZN(_3456_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8229_ (.A1(_3426_),
    .A2(_3425_),
    .B1(_3432_),
    .B2(_3433_),
    .C(_3456_),
    .ZN(_3457_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8230_ (.A1(_2782_),
    .A2(_3457_),
    .B(_3313_),
    .ZN(_3458_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8231_ (.A1(_3422_),
    .A2(_3425_),
    .B(_3458_),
    .ZN(_3459_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8232_ (.A1(_1314_),
    .A2(_3272_),
    .B(_3459_),
    .C(_3161_),
    .ZN(_0204_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8233_ (.A1(_2789_),
    .A2(_3423_),
    .ZN(_3460_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8234_ (.A1(_1321_),
    .A2(_3460_),
    .Z(_3461_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8235_ (.I(_3461_),
    .Z(_3462_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8236_ (.I(_2355_),
    .Z(_3463_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8237_ (.A1(_1657_),
    .A2(_4096_),
    .Z(_3464_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _8238_ (.A1(_1092_),
    .A2(_4111_),
    .Z(_3465_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _8239_ (.A1(_1092_),
    .A2(_4111_),
    .Z(_3466_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8240_ (.A1(_3465_),
    .A2(_3448_),
    .B(_3466_),
    .ZN(_3467_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8241_ (.A1(_3464_),
    .A2(_3467_),
    .ZN(_3468_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8242_ (.A1(_3464_),
    .A2(_3467_),
    .ZN(_3469_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8243_ (.A1(_3027_),
    .A2(_3469_),
    .ZN(_3470_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8244_ (.A1(_1674_),
    .A2(_3463_),
    .B1(_3468_),
    .B2(_3470_),
    .ZN(_3471_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8245_ (.A1(_3235_),
    .A2(_3471_),
    .B(_3455_),
    .ZN(_3472_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8246_ (.I(_3276_),
    .Z(_3473_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8247_ (.A1(_1321_),
    .A2(_3442_),
    .Z(_3474_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8248_ (.I(_0397_),
    .Z(_3475_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8249_ (.A1(_1321_),
    .A2(_0410_),
    .ZN(_3476_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8250_ (.A1(_1692_),
    .A2(_2869_),
    .B(_3476_),
    .ZN(_3477_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8251_ (.A1(_3475_),
    .A2(_3477_),
    .ZN(_3478_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8252_ (.A1(_1143_),
    .A2(_0463_),
    .B1(_3370_),
    .B2(_2382_),
    .C(_4360_),
    .ZN(_3479_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8253_ (.A1(_2531_),
    .A2(_3461_),
    .B(_3478_),
    .C(_3479_),
    .ZN(_3480_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8254_ (.A1(_3473_),
    .A2(_3474_),
    .B(_3480_),
    .ZN(_3481_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8255_ (.A1(_3282_),
    .A2(_3462_),
    .B1(_3481_),
    .B2(_3232_),
    .ZN(_3482_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8256_ (.A1(_3260_),
    .A2(_3462_),
    .ZN(_3483_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8257_ (.A1(_3175_),
    .A2(_3477_),
    .B(_3483_),
    .C(_3455_),
    .ZN(_3484_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8258_ (.A1(_3310_),
    .A2(_3484_),
    .ZN(_3485_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8259_ (.A1(_3472_),
    .A2(_3482_),
    .B(_3485_),
    .ZN(_3486_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8260_ (.I(_2497_),
    .Z(_3487_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _8261_ (.A1(\as2650.stack[3][6] ),
    .A2(_3302_),
    .B1(_3303_),
    .B2(\as2650.stack[2][6] ),
    .ZN(_3488_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _8262_ (.A1(\as2650.stack[1][6] ),
    .A2(_3242_),
    .B1(_3245_),
    .B2(\as2650.stack[0][6] ),
    .C(_0722_),
    .ZN(_3489_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _8263_ (.A1(\as2650.stack[5][6] ),
    .A2(_3241_),
    .B1(_3244_),
    .B2(\as2650.stack[4][6] ),
    .ZN(_3490_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _8264_ (.I(_3490_),
    .ZN(_3491_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _8265_ (.A1(\as2650.stack[7][6] ),
    .A2(_3250_),
    .B1(_3251_),
    .B2(\as2650.stack[6][6] ),
    .C(_3491_),
    .ZN(_3492_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _8266_ (.A1(_3488_),
    .A2(_3489_),
    .B1(_3492_),
    .B2(_1047_),
    .ZN(_3493_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8267_ (.A1(_3378_),
    .A2(_3462_),
    .ZN(_3494_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8268_ (.I(_3263_),
    .Z(_3495_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8269_ (.A1(_3487_),
    .A2(_3493_),
    .B(_3494_),
    .C(_3495_),
    .ZN(_3496_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _8270_ (.A1(_3273_),
    .A2(_3462_),
    .B1(_3486_),
    .B2(_3496_),
    .C(_3313_),
    .ZN(_3497_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8271_ (.A1(_1322_),
    .A2(_3269_),
    .B(_3497_),
    .ZN(_3498_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8272_ (.A1(_0335_),
    .A2(_3498_),
    .ZN(_0205_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8273_ (.I(_3391_),
    .Z(_3499_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8274_ (.A1(_1320_),
    .A2(_2788_),
    .A3(_3423_),
    .ZN(_3500_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8275_ (.A1(_1327_),
    .A2(_3500_),
    .Z(_3501_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8276_ (.I(_3501_),
    .Z(_3502_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _8277_ (.A1(\as2650.stack[3][7] ),
    .A2(_2389_),
    .B1(_1574_),
    .B2(\as2650.stack[2][7] ),
    .ZN(_3503_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _8278_ (.A1(\as2650.stack[1][7] ),
    .A2(_2456_),
    .B1(_3380_),
    .B2(\as2650.stack[0][7] ),
    .C(_1047_),
    .ZN(_3504_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _8279_ (.A1(\as2650.stack[5][7] ),
    .A2(_3242_),
    .B1(_3251_),
    .B2(\as2650.stack[6][7] ),
    .ZN(_3505_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _8280_ (.I(_3505_),
    .ZN(_3506_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _8281_ (.A1(\as2650.stack[7][7] ),
    .A2(_2389_),
    .B1(_3380_),
    .B2(\as2650.stack[4][7] ),
    .C(_3506_),
    .ZN(_3507_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _8282_ (.A1(_3503_),
    .A2(_3504_),
    .B1(_3507_),
    .B2(_0723_),
    .ZN(_3508_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8283_ (.A1(_2585_),
    .A2(_2884_),
    .ZN(_3509_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _8284_ (.A1(_1328_),
    .A2(_4415_),
    .B(_3509_),
    .C(_0813_),
    .ZN(_3510_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8285_ (.A1(_3194_),
    .A2(_3502_),
    .B(_3510_),
    .C(_0435_),
    .ZN(_3511_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8286_ (.I(_3281_),
    .Z(_3512_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _8287_ (.A1(_1320_),
    .A2(_3442_),
    .Z(_3513_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8288_ (.A1(_1328_),
    .A2(_3513_),
    .Z(_3514_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8289_ (.A1(_4262_),
    .A2(_4435_),
    .ZN(_3515_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8290_ (.A1(_2554_),
    .A2(_3293_),
    .B1(_3501_),
    .B2(_2595_),
    .ZN(_3516_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8291_ (.A1(_2536_),
    .A2(_3515_),
    .B(_3516_),
    .ZN(_3517_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8292_ (.A1(_3475_),
    .A2(_3510_),
    .B1(_3517_),
    .B2(_4048_),
    .ZN(_3518_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8293_ (.A1(_3441_),
    .A2(_3514_),
    .B(_3518_),
    .ZN(_3519_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8294_ (.A1(_2898_),
    .A2(_4096_),
    .B(_3469_),
    .ZN(_3520_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _8295_ (.A1(_2584_),
    .A2(_4073_),
    .A3(_3520_),
    .Z(_3521_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8296_ (.A1(_2552_),
    .A2(_3521_),
    .ZN(_3522_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8297_ (.A1(_0392_),
    .A2(_2723_),
    .B(_3234_),
    .C(_3522_),
    .ZN(_3523_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8298_ (.A1(_2712_),
    .A2(_3523_),
    .ZN(_3524_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8299_ (.A1(_3512_),
    .A2(_3502_),
    .B1(_3519_),
    .B2(_3238_),
    .C(_3524_),
    .ZN(_3525_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _8300_ (.A1(_2861_),
    .A2(_3511_),
    .A3(_3525_),
    .ZN(_3526_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8301_ (.A1(_3344_),
    .A2(_3502_),
    .B1(_3508_),
    .B2(_3258_),
    .C(_3526_),
    .ZN(_3527_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _8302_ (.A1(_2782_),
    .A2(_3527_),
    .Z(_3528_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8303_ (.A1(_3221_),
    .A2(_3502_),
    .B(_3271_),
    .ZN(_3529_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8304_ (.A1(_1328_),
    .A2(_3499_),
    .B1(_3528_),
    .B2(_3529_),
    .C(_0334_),
    .ZN(_0206_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8305_ (.A1(_1327_),
    .A2(_3500_),
    .ZN(_3530_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8306_ (.A1(_1379_),
    .A2(_3530_),
    .Z(_3531_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8307_ (.I(_3531_),
    .Z(_3532_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8308_ (.A1(_1379_),
    .A2(\as2650.pc[7] ),
    .A3(_3513_),
    .ZN(_3533_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8309_ (.A1(_2879_),
    .A2(_3513_),
    .B(_1380_),
    .ZN(_3534_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _8310_ (.A1(_4425_),
    .A2(_3473_),
    .A3(_3534_),
    .ZN(_3535_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8311_ (.A1(_3533_),
    .A2(_3535_),
    .ZN(_3536_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8312_ (.I(_3512_),
    .Z(_3537_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8313_ (.A1(_2584_),
    .A2(_4073_),
    .ZN(_3538_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8314_ (.A1(_0390_),
    .A2(_4073_),
    .ZN(_3539_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8315_ (.A1(_3538_),
    .A2(_3520_),
    .B(_3539_),
    .ZN(_3540_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8316_ (.A1(_2891_),
    .A2(_3540_),
    .ZN(_3541_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8317_ (.A1(_2362_),
    .A2(_3541_),
    .Z(_3542_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8318_ (.A1(_2361_),
    .A2(_2891_),
    .ZN(_3543_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8319_ (.A1(_2329_),
    .A2(_4436_),
    .B(_3543_),
    .ZN(_3544_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8320_ (.A1(_1380_),
    .A2(_2586_),
    .ZN(_3545_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8321_ (.A1(_0411_),
    .A2(_2955_),
    .B(_3545_),
    .C(_3475_),
    .ZN(_3546_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _8322_ (.A1(_2531_),
    .A2(_3531_),
    .B1(_3544_),
    .B2(_0358_),
    .C(_3546_),
    .ZN(_3547_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _8323_ (.A1(_4429_),
    .A2(_3542_),
    .B1(_3547_),
    .B2(_3139_),
    .ZN(_3548_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8324_ (.A1(_3537_),
    .A2(_3532_),
    .B1(_3548_),
    .B2(_3188_),
    .ZN(_3549_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8325_ (.A1(_0395_),
    .A2(_3536_),
    .A3(_3549_),
    .ZN(_3550_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8326_ (.I(_1511_),
    .Z(_3551_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _8327_ (.A1(_3487_),
    .A2(_0730_),
    .B1(_3551_),
    .B2(_3532_),
    .C(_3495_),
    .ZN(_3552_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8328_ (.A1(_1380_),
    .A2(_2538_),
    .ZN(_3553_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8329_ (.A1(_2385_),
    .A2(_2955_),
    .B(_3553_),
    .C(_1489_),
    .ZN(_3554_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8330_ (.I(_2712_),
    .Z(_3555_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8331_ (.A1(_3195_),
    .A2(_3532_),
    .B(_3554_),
    .C(_3555_),
    .ZN(_3556_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8332_ (.A1(_3552_),
    .A2(_3556_),
    .ZN(_3557_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8333_ (.A1(_3316_),
    .A2(_3532_),
    .B1(_3550_),
    .B2(_3557_),
    .C(_3220_),
    .ZN(_3558_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8334_ (.A1(_1381_),
    .A2(_3269_),
    .B(_3354_),
    .ZN(_3559_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8335_ (.A1(_3558_),
    .A2(_3559_),
    .ZN(_0207_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8336_ (.A1(_1379_),
    .A2(_3530_),
    .ZN(_3560_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8337_ (.A1(_1390_),
    .A2(_3560_),
    .Z(_3561_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8338_ (.I(_3561_),
    .Z(_3562_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _8339_ (.A1(_1389_),
    .A2(_3533_),
    .ZN(_3563_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _8340_ (.A1(_1390_),
    .A2(_3533_),
    .Z(_3564_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8341_ (.A1(_2965_),
    .A2(_0391_),
    .ZN(_3565_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8342_ (.A1(_0410_),
    .A2(_2984_),
    .B(_3565_),
    .ZN(_3566_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8343_ (.A1(_2366_),
    .A2(_2720_),
    .ZN(_3567_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8344_ (.A1(_3287_),
    .A2(_3567_),
    .B(_0357_),
    .ZN(_3568_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8345_ (.A1(_3475_),
    .A2(_3566_),
    .B1(_3561_),
    .B2(_2595_),
    .C(_3568_),
    .ZN(_3569_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _8346_ (.A1(_3441_),
    .A2(_3563_),
    .A3(_3564_),
    .B1(_3569_),
    .B2(_1488_),
    .ZN(_3570_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8347_ (.A1(_3238_),
    .A2(_3570_),
    .ZN(_3571_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8348_ (.A1(_2972_),
    .A2(_2720_),
    .A3(_3540_),
    .ZN(_3572_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8349_ (.A1(_2970_),
    .A2(_3572_),
    .Z(_3573_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8350_ (.A1(_3281_),
    .A2(_3562_),
    .B1(_3573_),
    .B2(_3234_),
    .C(_2548_),
    .ZN(_3574_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8351_ (.A1(_2728_),
    .A2(_3566_),
    .B1(_3562_),
    .B2(_0557_),
    .C(_4443_),
    .ZN(_3575_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8352_ (.A1(_3571_),
    .A2(_3574_),
    .B(_3575_),
    .ZN(_3576_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8353_ (.A1(_3433_),
    .A2(_0832_),
    .B1(_3426_),
    .B2(_3562_),
    .C(_3576_),
    .ZN(_3577_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8354_ (.A1(_2816_),
    .A2(_3577_),
    .B(_3313_),
    .ZN(_3578_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8355_ (.A1(_3422_),
    .A2(_3562_),
    .B(_3578_),
    .ZN(_3579_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8356_ (.A1(_1390_),
    .A2(_3499_),
    .B(_3579_),
    .C(_0349_),
    .ZN(_0208_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8357_ (.A1(\as2650.pc[9] ),
    .A2(_1378_),
    .A3(_3530_),
    .ZN(_3580_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8358_ (.A1(_1400_),
    .A2(_3580_),
    .Z(_3581_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8359_ (.I(_3581_),
    .Z(_3582_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8360_ (.A1(_3422_),
    .A2(_3582_),
    .ZN(_3583_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8361_ (.A1(_3000_),
    .A2(_0411_),
    .ZN(_3584_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8362_ (.A1(_1693_),
    .A2(_3024_),
    .B(_3584_),
    .ZN(_3585_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8363_ (.A1(_2370_),
    .A2(_2355_),
    .B(_4428_),
    .ZN(_3586_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8364_ (.A1(_2369_),
    .A2(_3027_),
    .B(_3586_),
    .ZN(_3587_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8365_ (.A1(_0399_),
    .A2(_3585_),
    .B1(_3581_),
    .B2(_2597_),
    .C(_3587_),
    .ZN(_3588_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _8366_ (.A1(_2972_),
    .A2(_2366_),
    .A3(_4435_),
    .A4(_3540_),
    .Z(_3589_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _8367_ (.A1(_2370_),
    .A2(_3589_),
    .Z(_3590_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8368_ (.A1(_2371_),
    .A2(_3589_),
    .B(_2354_),
    .ZN(_3591_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _8369_ (.A1(_4425_),
    .A2(_3588_),
    .B1(_3590_),
    .B2(_3591_),
    .ZN(_3592_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8370_ (.A1(_3188_),
    .A2(_3592_),
    .ZN(_3593_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8371_ (.A1(_3000_),
    .A2(_3563_),
    .Z(_3594_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8372_ (.A1(_3537_),
    .A2(_3582_),
    .B1(_3594_),
    .B2(_3278_),
    .C(_3033_),
    .ZN(_3595_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8373_ (.A1(_3593_),
    .A2(_3595_),
    .ZN(_3596_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8374_ (.A1(_3188_),
    .A2(_3585_),
    .ZN(_3597_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8375_ (.A1(_3339_),
    .A2(_3582_),
    .B(_3555_),
    .ZN(_3598_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _8376_ (.A1(_2497_),
    .A2(_0908_),
    .B1(_3551_),
    .B2(_3582_),
    .C(_3495_),
    .ZN(_3599_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8377_ (.A1(_3597_),
    .A2(_3598_),
    .B(_3599_),
    .ZN(_3600_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8378_ (.A1(_3596_),
    .A2(_3600_),
    .B(_3391_),
    .ZN(_3601_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8379_ (.A1(_1400_),
    .A2(_3499_),
    .B1(_3583_),
    .B2(_3601_),
    .C(_0334_),
    .ZN(_0209_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _8380_ (.A1(_1399_),
    .A2(_3580_),
    .ZN(_3602_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8381_ (.A1(_1407_),
    .A2(_3602_),
    .Z(_3603_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8382_ (.I(_3603_),
    .Z(_3604_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8383_ (.A1(_2903_),
    .A2(_3056_),
    .ZN(_3605_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8384_ (.A1(_1408_),
    .A2(_2538_),
    .B(_3605_),
    .C(_4049_),
    .ZN(_3606_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8385_ (.A1(_2713_),
    .A2(_3606_),
    .ZN(_3607_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8386_ (.A1(_2999_),
    .A2(_3563_),
    .ZN(_3608_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8387_ (.A1(_1408_),
    .A2(_3608_),
    .Z(_3609_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8388_ (.A1(_2374_),
    .A2(_2553_),
    .ZN(_3610_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _8389_ (.A1(_3367_),
    .A2(_3610_),
    .Z(_3611_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8390_ (.A1(_3436_),
    .A2(_3603_),
    .ZN(_3612_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _8391_ (.A1(_3473_),
    .A2(_3609_),
    .B1(_3611_),
    .B2(_3162_),
    .C(_3612_),
    .ZN(_3613_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8392_ (.A1(_3607_),
    .A2(_3613_),
    .B(_3232_),
    .ZN(_3614_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8393_ (.A1(_2374_),
    .A2(_3590_),
    .Z(_3615_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8394_ (.A1(_3537_),
    .A2(_3604_),
    .B1(_3615_),
    .B2(_3235_),
    .ZN(_3616_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8395_ (.A1(_0395_),
    .A2(_3614_),
    .A3(_3616_),
    .ZN(_3617_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8396_ (.A1(_3176_),
    .A2(_3604_),
    .B(_0436_),
    .ZN(_3618_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _8397_ (.A1(_3487_),
    .A2(_0978_),
    .B1(_3551_),
    .B2(_3604_),
    .C(_3495_),
    .ZN(_3619_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8398_ (.A1(_3606_),
    .A2(_3618_),
    .B(_3619_),
    .ZN(_3620_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8399_ (.A1(_3316_),
    .A2(_3604_),
    .B1(_3617_),
    .B2(_3620_),
    .C(_3220_),
    .ZN(_3621_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8400_ (.I(_3268_),
    .Z(_3622_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8401_ (.A1(_1409_),
    .A2(_3622_),
    .B(_3354_),
    .ZN(_3623_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8402_ (.A1(_3621_),
    .A2(_3623_),
    .ZN(_0210_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8403_ (.A1(_3069_),
    .A2(_3499_),
    .ZN(_3624_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8404_ (.A1(_1406_),
    .A2(_3602_),
    .ZN(_3625_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8405_ (.A1(_1416_),
    .A2(_3625_),
    .Z(_3626_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8406_ (.I(_3626_),
    .Z(_3627_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8407_ (.A1(\as2650.addr_buff[2] ),
    .A2(\as2650.addr_buff[3] ),
    .A3(_3589_),
    .ZN(_3628_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8408_ (.A1(_2378_),
    .A2(_3628_),
    .Z(_3629_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _8409_ (.I(_3401_),
    .ZN(_3630_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8410_ (.A1(_2378_),
    .A2(_2722_),
    .B(_3630_),
    .C(_3139_),
    .ZN(_3631_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8411_ (.A1(_4425_),
    .A2(_3629_),
    .B(_3631_),
    .C(_3162_),
    .ZN(_3632_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8412_ (.A1(_1406_),
    .A2(_2999_),
    .A3(_3563_),
    .ZN(_3633_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8413_ (.A1(_1416_),
    .A2(_3633_),
    .Z(_3634_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8414_ (.A1(_2384_),
    .A2(_3088_),
    .ZN(_3635_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8415_ (.A1(_3068_),
    .A2(_2537_),
    .B(_3635_),
    .ZN(_3636_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8416_ (.A1(_0425_),
    .A2(_3626_),
    .B(_1622_),
    .ZN(_3637_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8417_ (.A1(_0425_),
    .A2(_3636_),
    .B(_3637_),
    .ZN(_3638_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _8418_ (.A1(_3512_),
    .A2(_3627_),
    .B1(_3634_),
    .B2(_3277_),
    .C1(_3238_),
    .C2(_3638_),
    .ZN(_3639_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8419_ (.A1(_3555_),
    .A2(_3639_),
    .ZN(_3640_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8420_ (.A1(_3175_),
    .A2(_3627_),
    .ZN(_3641_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8421_ (.A1(_2473_),
    .A2(_3636_),
    .B(_3641_),
    .C(_3455_),
    .ZN(_3642_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8422_ (.A1(_3632_),
    .A2(_3640_),
    .B(_4368_),
    .C(_3642_),
    .ZN(_3643_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8423_ (.A1(_3433_),
    .A2(_1049_),
    .B1(_3344_),
    .B2(_3627_),
    .C(_2781_),
    .ZN(_3644_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8424_ (.A1(_3643_),
    .A2(_3644_),
    .ZN(_3645_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8425_ (.A1(_3273_),
    .A2(_3627_),
    .B(_3645_),
    .C(_3622_),
    .ZN(_3646_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8426_ (.I(_0469_),
    .Z(_3647_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8427_ (.A1(_3624_),
    .A2(_3646_),
    .B(_3647_),
    .ZN(_0211_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8428_ (.I(_0333_),
    .Z(_3648_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8429_ (.A1(_1422_),
    .A2(_3622_),
    .ZN(_3649_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8430_ (.I(\as2650.pc[13] ),
    .Z(_3650_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8431_ (.A1(_3068_),
    .A2(_1407_),
    .A3(_3602_),
    .ZN(_3651_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _8432_ (.A1(_3650_),
    .A2(_3651_),
    .ZN(_3652_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8433_ (.A1(_2597_),
    .A2(_3652_),
    .ZN(_3653_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _8434_ (.A1(_1422_),
    .A2(_0392_),
    .Z(_3654_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8435_ (.A1(_2380_),
    .A2(_0463_),
    .B1(_3654_),
    .B2(_0399_),
    .C(_4424_),
    .ZN(_3655_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8436_ (.A1(_2380_),
    .A2(_3463_),
    .B(_4429_),
    .ZN(_3656_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8437_ (.A1(_2374_),
    .A2(_2378_),
    .A3(_3590_),
    .ZN(_3657_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8438_ (.A1(_3653_),
    .A2(_3655_),
    .B1(_3656_),
    .B2(_3657_),
    .ZN(_3658_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8439_ (.A1(_3650_),
    .A2(_3651_),
    .Z(_3659_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8440_ (.A1(_1416_),
    .A2(_3633_),
    .ZN(_3660_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _8441_ (.A1(_3650_),
    .A2(_3660_),
    .ZN(_3661_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8442_ (.A1(_3512_),
    .A2(_3659_),
    .B1(_3661_),
    .B2(_3278_),
    .C(_3033_),
    .ZN(_3662_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8443_ (.A1(_3339_),
    .A2(_3658_),
    .B(_3662_),
    .ZN(_3663_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8444_ (.A1(_2472_),
    .A2(_3654_),
    .ZN(_3664_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8445_ (.A1(_3194_),
    .A2(_3659_),
    .B(_3664_),
    .C(_0435_),
    .ZN(_3665_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8446_ (.A1(_3433_),
    .A2(_1114_),
    .B1(_3426_),
    .B2(_3652_),
    .C(_3665_),
    .ZN(_3666_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8447_ (.A1(_3663_),
    .A2(_3666_),
    .B(_2816_),
    .ZN(_3667_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8448_ (.A1(_3422_),
    .A2(_3652_),
    .B(_3667_),
    .C(_3271_),
    .ZN(_3668_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _8449_ (.A1(_3648_),
    .A2(_3649_),
    .A3(_3668_),
    .ZN(_0212_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _8450_ (.A1(_3650_),
    .A2(_3068_),
    .A3(_1407_),
    .A4(_3602_),
    .ZN(_3669_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _8451_ (.A1(\as2650.pc[14] ),
    .A2(_3669_),
    .ZN(_3670_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8452_ (.A1(_1422_),
    .A2(_3660_),
    .ZN(_3671_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _8453_ (.A1(_1429_),
    .A2(_3473_),
    .A3(_3671_),
    .ZN(_3672_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _8454_ (.I(_3671_),
    .ZN(_3673_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8455_ (.A1(_3441_),
    .A2(_3673_),
    .B(_1756_),
    .ZN(_3674_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8456_ (.A1(\as2650.pc[14] ),
    .A2(_3674_),
    .ZN(_3675_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _8457_ (.A1(_0656_),
    .A2(_3463_),
    .A3(_3162_),
    .B(_3675_),
    .ZN(_3676_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8458_ (.A1(_3672_),
    .A2(_3676_),
    .B(_3232_),
    .ZN(_3677_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8459_ (.A1(_3537_),
    .A2(_3436_),
    .B(_3670_),
    .ZN(_3678_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8460_ (.A1(_2382_),
    .A2(_3463_),
    .A3(_3235_),
    .ZN(_3679_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _8461_ (.A1(_0395_),
    .A2(_3677_),
    .A3(_3678_),
    .A4(_3679_),
    .ZN(_3680_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _8462_ (.A1(_3487_),
    .A2(_1128_),
    .B1(_3551_),
    .B2(_3670_),
    .ZN(_3681_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8463_ (.A1(_1429_),
    .A2(_1755_),
    .B1(_3670_),
    .B2(_3339_),
    .C(_3555_),
    .ZN(_3682_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _8464_ (.A1(_2782_),
    .A2(_3681_),
    .A3(_3682_),
    .ZN(_3683_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8465_ (.A1(_3316_),
    .A2(_3670_),
    .B1(_3680_),
    .B2(_3683_),
    .C(_3271_),
    .ZN(_3684_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8466_ (.A1(_1429_),
    .A2(_3622_),
    .B(_3354_),
    .ZN(_3685_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8467_ (.A1(_3684_),
    .A2(_3685_),
    .ZN(_0213_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8468_ (.I(_4282_),
    .Z(_3686_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8469_ (.I(_3686_),
    .Z(_3687_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8470_ (.I(_2566_),
    .Z(_3688_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8471_ (.A1(_2762_),
    .A2(_0651_),
    .ZN(_3689_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8472_ (.A1(_3688_),
    .A2(_0660_),
    .B(_3689_),
    .ZN(_3690_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8473_ (.I(_3686_),
    .Z(_3691_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8474_ (.A1(_3691_),
    .A2(_0638_),
    .ZN(_3692_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8475_ (.I(_2943_),
    .Z(_3693_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8476_ (.A1(_3687_),
    .A2(_3690_),
    .B(_3692_),
    .C(_3693_),
    .ZN(_3694_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8477_ (.I(_1698_),
    .Z(_3695_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8478_ (.A1(_1541_),
    .A2(_3695_),
    .ZN(_3696_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8479_ (.A1(_1632_),
    .A2(_0368_),
    .A3(_1264_),
    .ZN(_3697_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8480_ (.I(_3697_),
    .Z(_3698_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8481_ (.A1(_0700_),
    .A2(_3698_),
    .ZN(_3699_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _8482_ (.A1(_0480_),
    .A2(_0491_),
    .A3(_0478_),
    .ZN(_3700_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8483_ (.I(_3700_),
    .Z(_3701_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8484_ (.A1(_0610_),
    .A2(_3701_),
    .B(_0574_),
    .ZN(_3702_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8485_ (.A1(_1923_),
    .A2(_1472_),
    .ZN(_3703_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8486_ (.A1(_3699_),
    .A2(_3702_),
    .B(_3703_),
    .C(_1700_),
    .ZN(_3704_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8487_ (.A1(_0489_),
    .A2(_3256_),
    .B(_3704_),
    .ZN(_3705_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _8488_ (.A1(_1695_),
    .A2(_1651_),
    .A3(_3705_),
    .ZN(_3706_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8489_ (.A1(_1752_),
    .A2(_1695_),
    .B1(_3696_),
    .B2(_3706_),
    .C(_4368_),
    .ZN(_3707_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8490_ (.A1(_2993_),
    .A2(_1839_),
    .B(_1691_),
    .ZN(_3708_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _8491_ (.A1(_4299_),
    .A2(_4315_),
    .A3(_4385_),
    .A4(_0572_),
    .ZN(_3709_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8492_ (.A1(_1493_),
    .A2(_4308_),
    .B1(_1763_),
    .B2(_4392_),
    .C(_3709_),
    .ZN(_3710_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8493_ (.A1(_3169_),
    .A2(_3710_),
    .ZN(_3711_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8494_ (.A1(_0420_),
    .A2(_2344_),
    .ZN(_3712_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8495_ (.A1(_1493_),
    .A2(_4314_),
    .B(_1531_),
    .ZN(_3713_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8496_ (.A1(_4057_),
    .A2(_0493_),
    .B(_4359_),
    .ZN(_3714_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8497_ (.A1(_1764_),
    .A2(_3714_),
    .B(_2341_),
    .ZN(_3715_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _8498_ (.A1(_2821_),
    .A2(_3712_),
    .A3(_3713_),
    .B(_3715_),
    .ZN(_3716_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _8499_ (.A1(_4400_),
    .A2(_4318_),
    .A3(_3343_),
    .A4(_1638_),
    .ZN(_3717_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8500_ (.A1(_2352_),
    .A2(_1512_),
    .ZN(_3718_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8501_ (.A1(_3168_),
    .A2(_1643_),
    .B(_0553_),
    .C(_1635_),
    .ZN(_3719_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8502_ (.A1(_4170_),
    .A2(_2343_),
    .B(_1630_),
    .C(_1248_),
    .ZN(_3720_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _8503_ (.A1(_0566_),
    .A2(_3718_),
    .A3(_3719_),
    .A4(_3720_),
    .ZN(_3721_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8504_ (.A1(_1493_),
    .A2(_0641_),
    .ZN(_3722_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8505_ (.A1(_4418_),
    .A2(_3722_),
    .B(_4335_),
    .ZN(_3723_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8506_ (.A1(_2344_),
    .A2(_3723_),
    .B(_1528_),
    .ZN(_3724_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _8507_ (.A1(_1642_),
    .A2(_3717_),
    .A3(_3721_),
    .A4(_3724_),
    .ZN(_3725_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _8508_ (.A1(_1628_),
    .A2(_3711_),
    .A3(_3716_),
    .A4(_3725_),
    .ZN(_3726_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8509_ (.I(_3726_),
    .Z(_3727_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _8510_ (.A1(_1534_),
    .A2(_1615_),
    .B1(_3707_),
    .B2(_3708_),
    .C(_3727_),
    .ZN(_3728_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8511_ (.A1(_3694_),
    .A2(_3728_),
    .ZN(_3729_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8512_ (.I(_3726_),
    .Z(_3730_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8513_ (.I(_3730_),
    .Z(_3731_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8514_ (.A1(_0698_),
    .A2(_3731_),
    .B(_2482_),
    .ZN(_3732_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8515_ (.A1(_3729_),
    .A2(_3732_),
    .ZN(_0214_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8516_ (.A1(_3688_),
    .A2(_0806_),
    .ZN(_3733_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8517_ (.I(_2693_),
    .Z(_3734_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8518_ (.A1(_3734_),
    .A2(_0802_),
    .B(_0354_),
    .ZN(_3735_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8519_ (.A1(_0355_),
    .A2(_0775_),
    .B1(_3733_),
    .B2(_3735_),
    .C(_3693_),
    .ZN(_3736_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8520_ (.A1(_2410_),
    .A2(_3308_),
    .ZN(_3737_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8521_ (.I(_3697_),
    .Z(_3738_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8522_ (.A1(\as2650.psl[1] ),
    .A2(_3698_),
    .ZN(_3739_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8523_ (.A1(_0702_),
    .A2(_3738_),
    .B(_0574_),
    .C(_3739_),
    .ZN(_3740_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8524_ (.A1(_1922_),
    .A2(_0503_),
    .B(_3740_),
    .ZN(_3741_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8525_ (.A1(_3737_),
    .A2(_3741_),
    .B(_1701_),
    .ZN(_3742_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _8526_ (.A1(_1534_),
    .A2(_1697_),
    .B1(_1698_),
    .B2(_0950_),
    .C(_1639_),
    .ZN(_3743_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _8527_ (.A1(_1677_),
    .A2(_1695_),
    .B1(_3742_),
    .B2(_3743_),
    .C(_3310_),
    .ZN(_3744_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8528_ (.A1(_4368_),
    .A2(_4218_),
    .ZN(_3745_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8529_ (.A1(_1691_),
    .A2(_3745_),
    .ZN(_3746_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _8530_ (.A1(_1541_),
    .A2(_1615_),
    .B1(_3744_),
    .B2(_3746_),
    .C(_3727_),
    .ZN(_3747_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8531_ (.A1(_3736_),
    .A2(_3747_),
    .ZN(_3748_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8532_ (.A1(_1540_),
    .A2(_3731_),
    .B(_2482_),
    .ZN(_3749_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8533_ (.A1(_3748_),
    .A2(_3749_),
    .ZN(_0215_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8534_ (.I(_3730_),
    .Z(_3750_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8535_ (.A1(_3734_),
    .A2(_0874_),
    .ZN(_3751_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8536_ (.A1(_3688_),
    .A2(_0896_),
    .B(_0354_),
    .ZN(_3752_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8537_ (.A1(_0355_),
    .A2(_1591_),
    .B1(_3751_),
    .B2(_3752_),
    .C(_3693_),
    .ZN(_3753_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8538_ (.I(_0454_),
    .Z(_3754_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8539_ (.I(_1640_),
    .Z(_3755_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8540_ (.A1(\as2650.overflow ),
    .A2(_3701_),
    .ZN(_3756_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8541_ (.A1(_1350_),
    .A2(_3698_),
    .B(_0573_),
    .ZN(_3757_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8542_ (.A1(_2005_),
    .A2(_0572_),
    .ZN(_3758_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8543_ (.A1(_3756_),
    .A2(_3757_),
    .B(_1700_),
    .C(_3758_),
    .ZN(_3759_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8544_ (.A1(_0815_),
    .A2(_3350_),
    .B(_3759_),
    .ZN(_3760_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8545_ (.A1(_1541_),
    .A2(_1697_),
    .B1(_1698_),
    .B2(_1550_),
    .C(_3760_),
    .ZN(_3761_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _8546_ (.A1(_1678_),
    .A2(_3754_),
    .B1(_3755_),
    .B2(_3761_),
    .C1(_0365_),
    .C2(_0791_),
    .ZN(_3762_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8547_ (.A1(_4214_),
    .A2(_0466_),
    .B(_3730_),
    .C(_3762_),
    .ZN(_3763_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _8548_ (.A1(_1545_),
    .A2(_3750_),
    .B1(_3753_),
    .B2(_3763_),
    .ZN(_3764_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8549_ (.A1(_3202_),
    .A2(_3764_),
    .ZN(_0216_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8550_ (.I(_2693_),
    .Z(_3765_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8551_ (.A1(_2929_),
    .A2(_0962_),
    .ZN(_3766_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8552_ (.A1(_3765_),
    .A2(_0948_),
    .B(_3766_),
    .C(_3686_),
    .ZN(_3767_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8553_ (.A1(_3691_),
    .A2(_0940_),
    .B(_3767_),
    .ZN(_3768_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8554_ (.A1(_1589_),
    .A2(_3768_),
    .ZN(_3769_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8555_ (.I(_1701_),
    .Z(_3770_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8556_ (.A1(\as2650.psu[3] ),
    .A2(_3738_),
    .ZN(_3771_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8557_ (.I(_3700_),
    .Z(_3772_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8558_ (.A1(_1212_),
    .A2(_3772_),
    .B(_2402_),
    .ZN(_3773_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8559_ (.A1(_1915_),
    .A2(_1472_),
    .B1(_3386_),
    .B2(_0489_),
    .ZN(_3774_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8560_ (.A1(_3771_),
    .A2(_3773_),
    .B(_3774_),
    .ZN(_3775_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8561_ (.A1(_3770_),
    .A2(_3775_),
    .ZN(_3776_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8562_ (.I(_1697_),
    .Z(_3777_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8563_ (.A1(_0791_),
    .A2(_3777_),
    .B1(_3695_),
    .B2(_2144_),
    .ZN(_3778_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8564_ (.A1(_3755_),
    .A2(_3776_),
    .A3(_3778_),
    .ZN(_3779_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _8565_ (.A1(_2373_),
    .A2(_3754_),
    .B1(_0426_),
    .B2(_1550_),
    .C1(_4212_),
    .C2(_2606_),
    .ZN(_3780_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8566_ (.A1(_3769_),
    .A2(_3779_),
    .A3(_3780_),
    .ZN(_3781_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8567_ (.A1(_0969_),
    .A2(_3750_),
    .B(_3038_),
    .ZN(_3782_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8568_ (.A1(_3731_),
    .A2(_3781_),
    .B(_3782_),
    .ZN(_0217_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8569_ (.A1(_1303_),
    .A2(_3727_),
    .ZN(_3783_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8570_ (.A1(_2762_),
    .A2(_1035_),
    .ZN(_3784_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8571_ (.A1(_3765_),
    .A2(_1015_),
    .B(_3686_),
    .ZN(_3785_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _8572_ (.A1(_3691_),
    .A2(_1009_),
    .B1(_3784_),
    .B2(_3785_),
    .ZN(_3786_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8573_ (.A1(_0555_),
    .A2(_3738_),
    .ZN(_3787_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8574_ (.A1(\as2650.psu[4] ),
    .A2(_3772_),
    .B(_1460_),
    .ZN(_3788_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8575_ (.A1(_2410_),
    .A2(_3415_),
    .ZN(_3789_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8576_ (.A1(_1865_),
    .A2(_0502_),
    .B(_1701_),
    .ZN(_3790_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _8577_ (.A1(_3787_),
    .A2(_3788_),
    .B(_3789_),
    .C(_3790_),
    .ZN(_3791_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _8578_ (.A1(_1550_),
    .A2(_1650_),
    .B1(_0793_),
    .B2(_1561_),
    .C(_1670_),
    .ZN(_3792_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _8579_ (.A1(_2376_),
    .A2(_1670_),
    .B1(_3791_),
    .B2(_3792_),
    .C(_0380_),
    .ZN(_3793_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8580_ (.A1(_4198_),
    .A2(_0438_),
    .B(_3726_),
    .C(_3793_),
    .ZN(_3794_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8581_ (.A1(_2144_),
    .A2(_0426_),
    .B1(_1589_),
    .B2(_3786_),
    .C(_3794_),
    .ZN(_3795_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _8582_ (.A1(_1508_),
    .A2(_3783_),
    .A3(_3795_),
    .ZN(_0218_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8583_ (.A1(_3734_),
    .A2(_1104_),
    .ZN(_3796_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8584_ (.A1(_3688_),
    .A2(_1086_),
    .B(_0354_),
    .ZN(_3797_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8585_ (.A1(_0355_),
    .A2(_1078_),
    .B1(_3796_),
    .B2(_3797_),
    .C(_3693_),
    .ZN(_3798_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _8586_ (.A1(\as2650.psu[5] ),
    .A2(_3700_),
    .Z(_3799_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8587_ (.A1(\as2650.psl[5] ),
    .A2(_3698_),
    .B(_1460_),
    .C(_3799_),
    .ZN(_3800_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _8588_ (.A1(_1864_),
    .A2(_0502_),
    .B1(_3432_),
    .B2(_0732_),
    .C(_1700_),
    .ZN(_3801_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8589_ (.A1(_2144_),
    .A2(_1696_),
    .B1(_0520_),
    .B2(_1668_),
    .ZN(_3802_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8590_ (.A1(_3800_),
    .A2(_3801_),
    .B(_3802_),
    .ZN(_3803_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8591_ (.A1(_1640_),
    .A2(_3803_),
    .ZN(_3804_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8592_ (.A1(_3726_),
    .A2(_3804_),
    .ZN(_3805_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8593_ (.A1(_1490_),
    .A2(_3754_),
    .B1(_0365_),
    .B2(_1028_),
    .C(_3805_),
    .ZN(_3806_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8594_ (.A1(_4204_),
    .A2(_0466_),
    .B(_3806_),
    .ZN(_3807_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8595_ (.A1(_3798_),
    .A2(_3807_),
    .ZN(_3808_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8596_ (.A1(_1312_),
    .A2(_3750_),
    .B(_2482_),
    .ZN(_3809_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8597_ (.A1(_3808_),
    .A2(_3809_),
    .ZN(_0219_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8598_ (.A1(_2762_),
    .A2(_1138_),
    .ZN(_3810_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8599_ (.A1(_3765_),
    .A2(_1154_),
    .B(_3691_),
    .ZN(_3811_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _8600_ (.A1(_3687_),
    .A2(_1177_),
    .B1(_3810_),
    .B2(_3811_),
    .C(_2814_),
    .ZN(_3812_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8601_ (.A1(_0815_),
    .A2(_3493_),
    .ZN(_3813_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _8602_ (.I(net28),
    .ZN(_3814_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8603_ (.A1(_1660_),
    .A2(_3701_),
    .ZN(_3815_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8604_ (.A1(_3814_),
    .A2(_3701_),
    .B(_3815_),
    .ZN(_3816_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8605_ (.A1(_4092_),
    .A2(_1472_),
    .B1(_2402_),
    .B2(_3816_),
    .ZN(_3817_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8606_ (.A1(_3813_),
    .A2(_3817_),
    .B(_0448_),
    .ZN(_3818_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8607_ (.A1(_1028_),
    .A2(_3777_),
    .B1(_3695_),
    .B2(_1619_),
    .C(_3818_),
    .ZN(_3819_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _8608_ (.A1(_1659_),
    .A2(_3754_),
    .B1(_3755_),
    .B2(_3819_),
    .C1(_0426_),
    .C2(_1090_),
    .ZN(_3820_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8609_ (.A1(_4188_),
    .A2(_0466_),
    .B(_3812_),
    .C(_3820_),
    .ZN(_3821_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8610_ (.A1(_1319_),
    .A2(_3750_),
    .B(_0351_),
    .ZN(_3822_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8611_ (.A1(_3731_),
    .A2(_3821_),
    .B(_3822_),
    .ZN(_0220_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8612_ (.A1(_3765_),
    .A2(_1228_),
    .ZN(_3823_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8613_ (.A1(_3734_),
    .A2(_1234_),
    .B(_3823_),
    .C(_3687_),
    .ZN(_3824_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8614_ (.A1(_3687_),
    .A2(_1209_),
    .B(_1589_),
    .C(_3824_),
    .ZN(_3825_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _8615_ (.A1(_1690_),
    .A2(_3738_),
    .Z(_3826_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8616_ (.A1(\as2650.psu[7] ),
    .A2(_3772_),
    .B(_1460_),
    .C(_3826_),
    .ZN(_3827_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _8617_ (.A1(_2230_),
    .A2(_0503_),
    .B1(_3508_),
    .B2(_0733_),
    .C(_3770_),
    .ZN(_3828_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8618_ (.A1(_3827_),
    .A2(_3828_),
    .B(_1699_),
    .ZN(_3829_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _8619_ (.A1(_2385_),
    .A2(_0678_),
    .B1(_1615_),
    .B2(_1139_),
    .C(_3730_),
    .ZN(_3830_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8620_ (.A1(_1217_),
    .A2(_2606_),
    .B1(_3755_),
    .B2(_3829_),
    .C(_3830_),
    .ZN(_3831_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8621_ (.A1(_1240_),
    .A2(_3727_),
    .B(_0351_),
    .ZN(_3832_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8622_ (.A1(_3825_),
    .A2(_3831_),
    .B(_3832_),
    .ZN(_0221_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _8623_ (.A1(_1346_),
    .A2(_1349_),
    .A3(_1351_),
    .A4(_1347_),
    .ZN(_3833_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8624_ (.I(_3833_),
    .Z(_3834_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8625_ (.I(_3833_),
    .Z(_3835_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8626_ (.A1(\as2650.stack[7][0] ),
    .A2(_3835_),
    .ZN(_3836_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8627_ (.A1(_2279_),
    .A2(_3834_),
    .B(_3836_),
    .ZN(_0222_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8628_ (.A1(\as2650.stack[7][1] ),
    .A2(_3835_),
    .ZN(_3837_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8629_ (.A1(_2285_),
    .A2(_3834_),
    .B(_3837_),
    .ZN(_0223_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8630_ (.A1(\as2650.stack[7][2] ),
    .A2(_3835_),
    .ZN(_3838_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8631_ (.A1(_2287_),
    .A2(_3834_),
    .B(_3838_),
    .ZN(_0224_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8632_ (.A1(\as2650.stack[7][3] ),
    .A2(_3835_),
    .ZN(_3839_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8633_ (.A1(_2289_),
    .A2(_3834_),
    .B(_3839_),
    .ZN(_0225_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8634_ (.I(_3833_),
    .Z(_3840_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8635_ (.I(_3833_),
    .Z(_3841_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8636_ (.A1(\as2650.stack[7][4] ),
    .A2(_3841_),
    .ZN(_3842_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8637_ (.A1(_2291_),
    .A2(_3840_),
    .B(_3842_),
    .ZN(_0226_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8638_ (.A1(\as2650.stack[7][5] ),
    .A2(_3841_),
    .ZN(_3843_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8639_ (.A1(_2295_),
    .A2(_3840_),
    .B(_3843_),
    .ZN(_0227_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8640_ (.A1(\as2650.stack[7][6] ),
    .A2(_3841_),
    .ZN(_3844_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8641_ (.A1(_2297_),
    .A2(_3840_),
    .B(_3844_),
    .ZN(_0228_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8642_ (.A1(\as2650.stack[7][7] ),
    .A2(_3841_),
    .ZN(_3845_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8643_ (.A1(_2299_),
    .A2(_3840_),
    .B(_3845_),
    .ZN(_0229_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _8644_ (.A1(_1436_),
    .A2(_1782_),
    .A3(_1783_),
    .ZN(_3846_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8645_ (.I(_3846_),
    .Z(_3847_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8646_ (.I(_3847_),
    .Z(_3848_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8647_ (.I(_3847_),
    .Z(_3849_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8648_ (.A1(\as2650.stack[7][8] ),
    .A2(_3849_),
    .ZN(_3850_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8649_ (.A1(_1781_),
    .A2(_3848_),
    .B(_3850_),
    .ZN(_0230_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8650_ (.I(_3846_),
    .Z(_3851_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8651_ (.A1(\as2650.stack[7][9] ),
    .A2(_3851_),
    .ZN(_3852_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8652_ (.A1(_1789_),
    .A2(_3848_),
    .B(_3852_),
    .ZN(_0231_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8653_ (.A1(\as2650.stack[7][10] ),
    .A2(_3851_),
    .ZN(_3853_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8654_ (.A1(_1792_),
    .A2(_3848_),
    .B(_3853_),
    .ZN(_0232_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8655_ (.A1(\as2650.stack[7][11] ),
    .A2(_3851_),
    .ZN(_3854_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8656_ (.A1(_1794_),
    .A2(_3848_),
    .B(_3854_),
    .ZN(_0233_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8657_ (.A1(\as2650.stack[7][12] ),
    .A2(_3851_),
    .ZN(_3855_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8658_ (.A1(_1796_),
    .A2(_3849_),
    .B(_3855_),
    .ZN(_0234_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8659_ (.A1(\as2650.stack[7][13] ),
    .A2(_3847_),
    .ZN(_3856_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8660_ (.A1(_1798_),
    .A2(_3849_),
    .B(_3856_),
    .ZN(_0235_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8661_ (.A1(\as2650.stack[7][14] ),
    .A2(_3847_),
    .ZN(_3857_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8662_ (.A1(_1800_),
    .A2(_3849_),
    .B(_3857_),
    .ZN(_0236_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _8663_ (.A1(_1436_),
    .A2(_1349_),
    .A3(_2280_),
    .A4(_1347_),
    .ZN(_3858_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8664_ (.I(_3858_),
    .Z(_3859_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8665_ (.I(_3858_),
    .Z(_3860_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8666_ (.A1(\as2650.stack[6][0] ),
    .A2(_3860_),
    .ZN(_3861_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8667_ (.A1(_2279_),
    .A2(_3859_),
    .B(_3861_),
    .ZN(_0237_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8668_ (.A1(\as2650.stack[6][1] ),
    .A2(_3860_),
    .ZN(_3862_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8669_ (.A1(_2285_),
    .A2(_3859_),
    .B(_3862_),
    .ZN(_0238_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8670_ (.A1(\as2650.stack[6][2] ),
    .A2(_3860_),
    .ZN(_3863_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8671_ (.A1(_2287_),
    .A2(_3859_),
    .B(_3863_),
    .ZN(_0239_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8672_ (.A1(\as2650.stack[6][3] ),
    .A2(_3860_),
    .ZN(_3864_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8673_ (.A1(_2289_),
    .A2(_3859_),
    .B(_3864_),
    .ZN(_0240_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8674_ (.I(_3858_),
    .Z(_3865_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8675_ (.I(_3858_),
    .Z(_3866_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8676_ (.A1(\as2650.stack[6][4] ),
    .A2(_3866_),
    .ZN(_3867_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8677_ (.A1(_2291_),
    .A2(_3865_),
    .B(_3867_),
    .ZN(_0241_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8678_ (.A1(\as2650.stack[6][5] ),
    .A2(_3866_),
    .ZN(_3868_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8679_ (.A1(_2295_),
    .A2(_3865_),
    .B(_3868_),
    .ZN(_0242_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8680_ (.A1(\as2650.stack[6][6] ),
    .A2(_3866_),
    .ZN(_3869_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8681_ (.A1(_2297_),
    .A2(_3865_),
    .B(_3869_),
    .ZN(_0243_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8682_ (.A1(\as2650.stack[6][7] ),
    .A2(_3866_),
    .ZN(_3870_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8683_ (.A1(_2299_),
    .A2(_3865_),
    .B(_3870_),
    .ZN(_0244_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _8684_ (.A1(_1243_),
    .A2(_3380_),
    .A3(_1782_),
    .ZN(_3871_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8685_ (.I(_3871_),
    .Z(_3872_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8686_ (.I(_3872_),
    .Z(_3873_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8687_ (.I(_3872_),
    .Z(_3874_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8688_ (.A1(\as2650.stack[5][8] ),
    .A2(_3874_),
    .ZN(_3875_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8689_ (.A1(_1781_),
    .A2(_3873_),
    .B(_3875_),
    .ZN(_0245_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8690_ (.I(_3871_),
    .Z(_3876_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8691_ (.A1(\as2650.stack[5][9] ),
    .A2(_3876_),
    .ZN(_3877_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8692_ (.A1(_1789_),
    .A2(_3873_),
    .B(_3877_),
    .ZN(_0246_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8693_ (.A1(\as2650.stack[5][10] ),
    .A2(_3876_),
    .ZN(_3878_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8694_ (.A1(_1792_),
    .A2(_3873_),
    .B(_3878_),
    .ZN(_0247_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8695_ (.A1(\as2650.stack[5][11] ),
    .A2(_3876_),
    .ZN(_3879_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8696_ (.A1(_1794_),
    .A2(_3873_),
    .B(_3879_),
    .ZN(_0248_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8697_ (.A1(\as2650.stack[5][12] ),
    .A2(_3876_),
    .ZN(_3880_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8698_ (.A1(_1796_),
    .A2(_3874_),
    .B(_3880_),
    .ZN(_0249_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8699_ (.A1(\as2650.stack[5][13] ),
    .A2(_3872_),
    .ZN(_3881_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8700_ (.A1(_1798_),
    .A2(_3874_),
    .B(_3881_),
    .ZN(_0250_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8701_ (.A1(\as2650.stack[5][14] ),
    .A2(_3872_),
    .ZN(_3882_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8702_ (.A1(_1800_),
    .A2(_3874_),
    .B(_3882_),
    .ZN(_0251_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8703_ (.A1(_1633_),
    .A2(_1132_),
    .ZN(_3883_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8704_ (.I(_0741_),
    .Z(_3884_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8705_ (.I(_3884_),
    .Z(_3885_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8706_ (.A1(_0480_),
    .A2(_0570_),
    .ZN(_3886_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _8707_ (.A1(_0468_),
    .A2(_3884_),
    .A3(_3886_),
    .ZN(_3887_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8708_ (.I(_3887_),
    .Z(_3888_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8709_ (.A1(_3885_),
    .A2(_1924_),
    .B1(_3888_),
    .B2(\as2650.r123[1][0] ),
    .ZN(_3889_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8710_ (.A1(_0696_),
    .A2(_3883_),
    .B(_3889_),
    .ZN(_0252_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8711_ (.I(_3887_),
    .Z(_3890_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8712_ (.A1(\as2650.r123[1][1] ),
    .A2(_3890_),
    .ZN(_3891_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8713_ (.I(_3884_),
    .Z(_3892_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8714_ (.I(_3886_),
    .Z(_3893_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8715_ (.A1(_3892_),
    .A2(_2309_),
    .B1(_3893_),
    .B2(_0811_),
    .ZN(_3894_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8716_ (.A1(_3891_),
    .A2(_3894_),
    .ZN(_0253_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8717_ (.A1(\as2650.r123[1][2] ),
    .A2(_3890_),
    .ZN(_3895_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8718_ (.A1(_3892_),
    .A2(_2312_),
    .B1(_3893_),
    .B2(_0901_),
    .ZN(_3896_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8719_ (.A1(_3895_),
    .A2(_3896_),
    .ZN(_0254_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8720_ (.A1(_3885_),
    .A2(_2314_),
    .B1(_3888_),
    .B2(\as2650.r123[1][3] ),
    .ZN(_3897_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8721_ (.A1(_0967_),
    .A2(_3883_),
    .B(_3897_),
    .ZN(_0255_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8722_ (.A1(\as2650.r123[1][4] ),
    .A2(_3890_),
    .ZN(_3898_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8723_ (.A1(_3892_),
    .A2(_2317_),
    .B1(_3893_),
    .B2(_1039_),
    .ZN(_3899_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8724_ (.A1(_3898_),
    .A2(_3899_),
    .ZN(_0256_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8725_ (.I(_0741_),
    .Z(_3900_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8726_ (.I(_3900_),
    .Z(_3901_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8727_ (.A1(_3901_),
    .A2(_2320_),
    .ZN(_3902_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8728_ (.A1(_1108_),
    .A2(_3893_),
    .B1(_3890_),
    .B2(\as2650.r123[1][5] ),
    .ZN(_3903_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8729_ (.A1(_3902_),
    .A2(_3903_),
    .ZN(_0257_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8730_ (.A1(_3885_),
    .A2(_2324_),
    .B1(_3888_),
    .B2(\as2650.r123[1][6] ),
    .ZN(_3904_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8731_ (.A1(_1179_),
    .A2(_3883_),
    .B(_3904_),
    .ZN(_0258_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8732_ (.A1(_3885_),
    .A2(_2326_),
    .B1(_3888_),
    .B2(\as2650.r123[1][7] ),
    .ZN(_3905_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8733_ (.A1(_1238_),
    .A2(_3883_),
    .B(_3905_),
    .ZN(_0259_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8734_ (.A1(_1729_),
    .A2(_1132_),
    .ZN(_3906_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8735_ (.A1(_1466_),
    .A2(_0570_),
    .ZN(_3907_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _8736_ (.A1(_0468_),
    .A2(_3884_),
    .A3(_3907_),
    .ZN(_3908_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8737_ (.I(_3908_),
    .Z(_3909_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8738_ (.A1(_3900_),
    .A2(_2036_),
    .B1(_3909_),
    .B2(\as2650.r123[2][0] ),
    .ZN(_3910_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8739_ (.A1(_0696_),
    .A2(_3906_),
    .B(_3910_),
    .ZN(_0260_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8740_ (.I(_3907_),
    .Z(_3911_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8741_ (.I(_3908_),
    .Z(_3912_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8742_ (.A1(_0811_),
    .A2(_3911_),
    .B1(_3912_),
    .B2(\as2650.r123[2][1] ),
    .ZN(_3913_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8743_ (.A1(_3901_),
    .A2(_2094_),
    .ZN(_3914_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8744_ (.A1(_3913_),
    .A2(_3914_),
    .ZN(_0261_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8745_ (.A1(_0901_),
    .A2(_3911_),
    .B1(_3912_),
    .B2(\as2650.r123[2][2] ),
    .ZN(_3915_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8746_ (.A1(_3901_),
    .A2(_2141_),
    .ZN(_3916_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8747_ (.A1(_3915_),
    .A2(_3916_),
    .ZN(_0262_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8748_ (.A1(_3900_),
    .A2(_2177_),
    .B1(_3909_),
    .B2(\as2650.r123[2][3] ),
    .ZN(_3917_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8749_ (.A1(_0967_),
    .A2(_3906_),
    .B(_3917_),
    .ZN(_0263_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8750_ (.A1(_1039_),
    .A2(_3911_),
    .B1(_3909_),
    .B2(\as2650.r123[2][4] ),
    .ZN(_3918_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _8751_ (.A1(_0551_),
    .A2(_0740_),
    .A3(_2198_),
    .B(_3918_),
    .ZN(_0264_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8752_ (.A1(_1108_),
    .A2(_3911_),
    .B1(_3912_),
    .B2(\as2650.r123[2][5] ),
    .ZN(_3919_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8753_ (.A1(_3901_),
    .A2(_2236_),
    .ZN(_3920_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8754_ (.A1(_3919_),
    .A2(_3920_),
    .ZN(_0265_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8755_ (.A1(_3900_),
    .A2(_2261_),
    .B1(_3909_),
    .B2(\as2650.r123[2][6] ),
    .ZN(_3921_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8756_ (.A1(_1179_),
    .A2(_3906_),
    .B(_3921_),
    .ZN(_0266_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8757_ (.A1(\as2650.r123[2][7] ),
    .A2(_3912_),
    .ZN(_3922_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8758_ (.A1(_3892_),
    .A2(_2276_),
    .ZN(_3923_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8759_ (.A1(_1238_),
    .A2(_3906_),
    .B(_3922_),
    .C(_3923_),
    .ZN(_0267_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8760_ (.A1(_2280_),
    .A2(_0715_),
    .A3(_1270_),
    .ZN(_3924_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8761_ (.I(_3924_),
    .Z(_3925_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8762_ (.I(_3924_),
    .Z(_3926_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8763_ (.A1(\as2650.stack[4][0] ),
    .A2(_3926_),
    .ZN(_3927_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8764_ (.A1(_2279_),
    .A2(_3925_),
    .B(_3927_),
    .ZN(_0268_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8765_ (.A1(\as2650.stack[4][1] ),
    .A2(_3926_),
    .ZN(_3928_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8766_ (.A1(_2285_),
    .A2(_3925_),
    .B(_3928_),
    .ZN(_0269_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8767_ (.A1(\as2650.stack[4][2] ),
    .A2(_3926_),
    .ZN(_3929_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8768_ (.A1(_2287_),
    .A2(_3925_),
    .B(_3929_),
    .ZN(_0270_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8769_ (.A1(\as2650.stack[4][3] ),
    .A2(_3926_),
    .ZN(_3930_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8770_ (.A1(_2289_),
    .A2(_3925_),
    .B(_3930_),
    .ZN(_0271_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8771_ (.I(_3924_),
    .Z(_3931_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8772_ (.I(_3924_),
    .Z(_3932_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8773_ (.A1(\as2650.stack[4][4] ),
    .A2(_3932_),
    .ZN(_3933_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8774_ (.A1(_2291_),
    .A2(_3931_),
    .B(_3933_),
    .ZN(_0272_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8775_ (.A1(\as2650.stack[4][5] ),
    .A2(_3932_),
    .ZN(_3934_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8776_ (.A1(_2295_),
    .A2(_3931_),
    .B(_3934_),
    .ZN(_0273_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8777_ (.A1(\as2650.stack[4][6] ),
    .A2(_3932_),
    .ZN(_3935_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8778_ (.A1(_2297_),
    .A2(_3931_),
    .B(_3935_),
    .ZN(_0274_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8779_ (.A1(\as2650.stack[4][7] ),
    .A2(_3932_),
    .ZN(_3936_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8780_ (.A1(_2299_),
    .A2(_3931_),
    .B(_3936_),
    .ZN(_0275_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8781_ (.A1(_1680_),
    .A2(_1754_),
    .ZN(_3937_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8782_ (.A1(_2993_),
    .A2(_1761_),
    .B(_3937_),
    .ZN(_0276_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8783_ (.A1(_2377_),
    .A2(_1754_),
    .ZN(_3938_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8784_ (.A1(_0321_),
    .A2(_1761_),
    .B(_3938_),
    .ZN(_0277_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8785_ (.I(_3378_),
    .Z(_3939_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8786_ (.A1(_1479_),
    .A2(_2639_),
    .ZN(_3940_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _8787_ (.A1(_0460_),
    .A2(_2336_),
    .A3(_0389_),
    .B1(_0360_),
    .B2(_0490_),
    .ZN(_3941_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _8788_ (.A1(_4424_),
    .A2(_3515_),
    .B1(_3941_),
    .B2(_4436_),
    .C(_4301_),
    .ZN(_3942_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8789_ (.A1(_0383_),
    .A2(_0442_),
    .B(_3370_),
    .C(_0388_),
    .ZN(_3943_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8790_ (.A1(_2471_),
    .A2(_0388_),
    .B(_2336_),
    .ZN(_3944_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8791_ (.A1(_0449_),
    .A2(_1471_),
    .B(_0428_),
    .C(_0677_),
    .ZN(_3945_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8792_ (.A1(_3943_),
    .A2(_3944_),
    .B(_3945_),
    .ZN(_3946_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8793_ (.A1(_4235_),
    .A2(_1258_),
    .B(_1478_),
    .C(_0429_),
    .ZN(_3947_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _8794_ (.A1(_4423_),
    .A2(_1249_),
    .B1(_1756_),
    .B2(_1258_),
    .ZN(_3948_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8795_ (.A1(_4367_),
    .A2(_3948_),
    .ZN(_3949_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8796_ (.A1(_3947_),
    .A2(_3949_),
    .ZN(_3950_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8797_ (.A1(_3168_),
    .A2(_0739_),
    .ZN(_3951_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8798_ (.A1(_4248_),
    .A2(_0368_),
    .A3(_1264_),
    .ZN(_3952_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _8799_ (.A1(_3952_),
    .A2(_0502_),
    .A3(_1248_),
    .A4(_1476_),
    .ZN(_3953_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8800_ (.A1(_3700_),
    .A2(_3951_),
    .B(_3953_),
    .C(_4308_),
    .ZN(_3954_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8801_ (.A1(_1630_),
    .A2(_3954_),
    .ZN(_3955_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _8802_ (.A1(_3133_),
    .A2(_3946_),
    .A3(_3950_),
    .A4(_3955_),
    .ZN(_3956_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _8803_ (.A1(_0423_),
    .A2(_1462_),
    .B1(_3942_),
    .B2(_3194_),
    .C(_3956_),
    .ZN(_3957_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8804_ (.A1(_3939_),
    .A2(_3940_),
    .B(_3957_),
    .ZN(_3958_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8805_ (.I(_1643_),
    .Z(_3959_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8806_ (.A1(_1350_),
    .A2(_1574_),
    .Z(_3960_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8807_ (.A1(_0877_),
    .A2(_3959_),
    .ZN(_3961_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8808_ (.A1(_3959_),
    .A2(_3960_),
    .B(_3961_),
    .C(_0733_),
    .ZN(_3962_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8809_ (.A1(_0733_),
    .A2(_0973_),
    .B(_3962_),
    .C(_3195_),
    .ZN(_3963_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8810_ (.A1(_1497_),
    .A2(_3181_),
    .B(_3963_),
    .C(_3939_),
    .ZN(_3964_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8811_ (.A1(_3258_),
    .A2(_0723_),
    .B1(_3960_),
    .B2(_0424_),
    .ZN(_3965_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8812_ (.A1(_3964_),
    .A2(_3965_),
    .ZN(_3966_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8813_ (.A1(_2280_),
    .A2(_3958_),
    .B(_0351_),
    .ZN(_3967_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8814_ (.A1(_3958_),
    .A2(_3966_),
    .B(_3967_),
    .ZN(_0278_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8815_ (.A1(_3250_),
    .A2(_3303_),
    .ZN(_3968_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8816_ (.A1(_3959_),
    .A2(_3968_),
    .B(_0732_),
    .ZN(_3969_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8817_ (.A1(_0778_),
    .A2(_3959_),
    .B(_3969_),
    .ZN(_3970_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8818_ (.A1(_2410_),
    .A2(_3968_),
    .B(_4361_),
    .ZN(_3971_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _8819_ (.A1(_1463_),
    .A2(_2365_),
    .A3(_1496_),
    .B1(_3970_),
    .B2(_3971_),
    .ZN(_3972_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8820_ (.A1(_1510_),
    .A2(_3972_),
    .ZN(_3973_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8821_ (.A1(_1477_),
    .A2(_3968_),
    .B(_3310_),
    .ZN(_3974_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8822_ (.A1(_0424_),
    .A2(_3968_),
    .B1(_3973_),
    .B2(_3974_),
    .ZN(_3975_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8823_ (.A1(_1499_),
    .A2(_1677_),
    .ZN(_3976_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8824_ (.A1(_3426_),
    .A2(_3976_),
    .B(_3957_),
    .ZN(_3977_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8825_ (.I0(_1349_),
    .I1(_3975_),
    .S(_3977_),
    .Z(_3978_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _8826_ (.A1(_1689_),
    .A2(_3978_),
    .Z(_3979_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8827_ (.I(_3979_),
    .Z(_0279_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8828_ (.A1(_2473_),
    .A2(_1752_),
    .ZN(_3980_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8829_ (.A1(_3344_),
    .A2(_3980_),
    .B(_3957_),
    .ZN(_3981_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8830_ (.A1(_3176_),
    .A2(_1644_),
    .ZN(_3982_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8831_ (.A1(_3982_),
    .A2(_3939_),
    .ZN(_3983_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _8832_ (.A1(_1644_),
    .A2(_3167_),
    .B1(_3171_),
    .B2(_1497_),
    .ZN(_3984_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8833_ (.A1(_1436_),
    .A2(_3983_),
    .B1(_3984_),
    .B2(_3939_),
    .ZN(_3985_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8834_ (.A1(_1346_),
    .A2(_3981_),
    .ZN(_3986_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8835_ (.A1(_3981_),
    .A2(_3985_),
    .B(_3986_),
    .C(_0349_),
    .ZN(_0280_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8836_ (.A1(_1614_),
    .A2(_3777_),
    .ZN(_3987_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8837_ (.A1(_4251_),
    .A2(_2343_),
    .ZN(_3988_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _8838_ (.A1(_0454_),
    .A2(_0364_),
    .A3(_1515_),
    .A4(_3988_),
    .ZN(_3989_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _8839_ (.A1(_1625_),
    .A2(_1641_),
    .A3(_1634_),
    .A4(_3989_),
    .ZN(_3990_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _8840_ (.I(_3990_),
    .ZN(_3991_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8841_ (.A1(_3169_),
    .A2(_3952_),
    .B(_0574_),
    .C(_1636_),
    .ZN(_3992_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8842_ (.A1(_1212_),
    .A2(_2472_),
    .B(_1626_),
    .ZN(_3993_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _8843_ (.A1(_3772_),
    .A2(_0479_),
    .A3(_3992_),
    .A4(_3993_),
    .ZN(_3994_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8844_ (.A1(_1630_),
    .A2(_3991_),
    .A3(_3994_),
    .ZN(_3995_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8845_ (.A1(_3987_),
    .A2(_3980_),
    .B(_3995_),
    .ZN(_3996_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8846_ (.A1(_1732_),
    .A2(_3171_),
    .B(_3167_),
    .C(_3770_),
    .ZN(_3997_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8847_ (.A1(_1139_),
    .A2(_3777_),
    .B1(_3695_),
    .B2(_1534_),
    .C(_1614_),
    .ZN(_3998_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8848_ (.A1(_3997_),
    .A2(_3998_),
    .ZN(_3999_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8849_ (.A1(_3996_),
    .A2(_3999_),
    .ZN(_4000_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8850_ (.A1(_0925_),
    .A2(_0934_),
    .ZN(_4001_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8851_ (.A1(_4001_),
    .A2(_0997_),
    .ZN(_4002_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8852_ (.A1(_4002_),
    .A2(_1596_),
    .B(_1606_),
    .ZN(_4003_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8853_ (.A1(_1192_),
    .A2(_1196_),
    .B(_1200_),
    .C(_1004_),
    .ZN(_4004_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8854_ (.A1(_0931_),
    .A2(_4003_),
    .B(_4004_),
    .ZN(_4005_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _8855_ (.A1(_2961_),
    .A2(_0914_),
    .A3(_4005_),
    .ZN(_4006_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _8856_ (.A1(_0610_),
    .A2(_3996_),
    .B1(_4000_),
    .B2(_4006_),
    .ZN(_4007_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8857_ (.A1(_3202_),
    .A2(_4007_),
    .ZN(_0281_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8858_ (.A1(_1491_),
    .A2(_3987_),
    .B(_3995_),
    .ZN(_4008_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8859_ (.A1(_3195_),
    .A2(_1476_),
    .B(_1503_),
    .C(_3770_),
    .ZN(_4009_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8860_ (.A1(_3802_),
    .A2(_4009_),
    .ZN(_4010_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _8861_ (.A1(_0931_),
    .A2(_0996_),
    .A3(_1008_),
    .ZN(_4011_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8862_ (.A1(_0306_),
    .A2(_4011_),
    .ZN(_4012_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8863_ (.A1(_0387_),
    .A2(_4010_),
    .B(_4012_),
    .ZN(_4013_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8864_ (.A1(\as2650.psl[5] ),
    .A2(_4008_),
    .ZN(_4014_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8865_ (.A1(_4008_),
    .A2(_4013_),
    .B(_4014_),
    .C(_0349_),
    .ZN(_0282_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8866_ (.A1(_0489_),
    .A2(_3951_),
    .B1(_3940_),
    .B2(_4402_),
    .ZN(_4015_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8867_ (.A1(_1626_),
    .A2(_4015_),
    .ZN(_4016_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _8868_ (.A1(_0485_),
    .A2(_1631_),
    .A3(_3990_),
    .A4(_4016_),
    .ZN(_4017_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8869_ (.I0(_1192_),
    .I1(_1193_),
    .S(_1208_),
    .Z(_4018_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8870_ (.A1(_1732_),
    .A2(_3180_),
    .ZN(_4019_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8871_ (.A1(_1691_),
    .A2(_3182_),
    .A3(_4019_),
    .ZN(_4020_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8872_ (.A1(_0387_),
    .A2(_4018_),
    .B(_4017_),
    .C(_4020_),
    .ZN(_4021_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8873_ (.A1(\as2650.overflow ),
    .A2(_4017_),
    .B(_4021_),
    .ZN(_4022_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8874_ (.A1(_3202_),
    .A2(_4022_),
    .ZN(_0283_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8875_ (.A1(_3174_),
    .A2(_2377_),
    .ZN(_4023_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8876_ (.A1(_0486_),
    .A2(_1461_),
    .ZN(_4024_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _8877_ (.A1(_0432_),
    .A2(_1509_),
    .A3(_2498_),
    .A4(_2989_),
    .ZN(_4025_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8878_ (.A1(_0480_),
    .A2(_3208_),
    .A3(_4025_),
    .ZN(_4026_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8879_ (.A1(_1622_),
    .A2(_1495_),
    .B(_4026_),
    .ZN(_4027_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _8880_ (.A1(_1464_),
    .A2(_1475_),
    .A3(_4024_),
    .A4(_4027_),
    .ZN(_4028_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8881_ (.A1(_4023_),
    .A2(_4028_),
    .B(_0555_),
    .ZN(_4029_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8882_ (.A1(_1732_),
    .A2(_3190_),
    .B(_4028_),
    .ZN(_4030_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8883_ (.A1(_3191_),
    .A2(_4030_),
    .ZN(_4031_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8884_ (.A1(_4029_),
    .A2(_4031_),
    .B(_3647_),
    .ZN(_0284_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8885_ (.A1(_3184_),
    .A2(_4028_),
    .B(_1212_),
    .ZN(_4032_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8886_ (.A1(_3185_),
    .A2(_4030_),
    .ZN(_4033_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8887_ (.A1(_4032_),
    .A2(_4033_),
    .B(_3647_),
    .ZN(_0285_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8888_ (.A1(_3976_),
    .A2(_4028_),
    .B(\as2650.psl[1] ),
    .ZN(_4034_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8889_ (.A1(_3178_),
    .A2(_4030_),
    .ZN(_4035_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8890_ (.A1(_4034_),
    .A2(_4035_),
    .B(_3647_),
    .ZN(_0286_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8891_ (.A1(_0494_),
    .A2(_0666_),
    .B(_4398_),
    .C(_4025_),
    .ZN(_4036_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _8892_ (.A1(_1654_),
    .A2(_1461_),
    .A3(_1470_),
    .A4(_4036_),
    .Z(_4037_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8893_ (.A1(_3196_),
    .A2(_4037_),
    .B(net28),
    .ZN(_4038_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8894_ (.A1(_4051_),
    .A2(_1497_),
    .B(_4037_),
    .ZN(_4039_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8895_ (.A1(_3197_),
    .A2(_4039_),
    .ZN(_4040_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8896_ (.A1(_4038_),
    .A2(_4040_),
    .B(_3648_),
    .ZN(_0287_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8897_ (.A1(_4023_),
    .A2(_4037_),
    .B(\as2650.psu[4] ),
    .ZN(_4041_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8898_ (.A1(_3191_),
    .A2(_4039_),
    .ZN(_4042_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8899_ (.A1(_4041_),
    .A2(_4042_),
    .B(_3648_),
    .ZN(_0288_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8900_ (.A1(_3184_),
    .A2(_4037_),
    .B(\as2650.psu[3] ),
    .ZN(_4043_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8901_ (.A1(_3185_),
    .A2(_4039_),
    .ZN(_4044_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8902_ (.A1(_4043_),
    .A2(_4044_),
    .B(_3648_),
    .ZN(_0289_));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8903_ (.D(_0014_),
    .CLK(clknet_leaf_63_wb_clk_i),
    .Q(\as2650.r123[3][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8904_ (.D(_0015_),
    .CLK(clknet_leaf_76_wb_clk_i),
    .Q(\as2650.r123[3][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8905_ (.D(_0016_),
    .CLK(clknet_leaf_60_wb_clk_i),
    .Q(\as2650.r123[3][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8906_ (.D(_0017_),
    .CLK(clknet_leaf_60_wb_clk_i),
    .Q(\as2650.r123[3][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8907_ (.D(_0018_),
    .CLK(clknet_leaf_63_wb_clk_i),
    .Q(\as2650.r123[3][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8908_ (.D(_0019_),
    .CLK(clknet_leaf_66_wb_clk_i),
    .Q(\as2650.r123[3][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8909_ (.D(_0020_),
    .CLK(clknet_leaf_75_wb_clk_i),
    .Q(\as2650.r123[3][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8910_ (.D(_0021_),
    .CLK(clknet_leaf_76_wb_clk_i),
    .Q(\as2650.r123[3][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8911_ (.D(_0022_),
    .CLK(clknet_leaf_68_wb_clk_i),
    .Q(\as2650.r123[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8912_ (.D(_0023_),
    .CLK(clknet_leaf_68_wb_clk_i),
    .Q(\as2650.r123[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8913_ (.D(_0024_),
    .CLK(clknet_leaf_68_wb_clk_i),
    .Q(\as2650.r123[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8914_ (.D(_0025_),
    .CLK(clknet_leaf_68_wb_clk_i),
    .Q(\as2650.r123[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8915_ (.D(_0026_),
    .CLK(clknet_leaf_68_wb_clk_i),
    .Q(\as2650.r123[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8916_ (.D(_0027_),
    .CLK(clknet_leaf_68_wb_clk_i),
    .Q(\as2650.r123[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8917_ (.D(_0028_),
    .CLK(clknet_leaf_68_wb_clk_i),
    .Q(\as2650.r123[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8918_ (.D(_0029_),
    .CLK(clknet_3_1__leaf_wb_clk_i),
    .Q(\as2650.r123[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8919_ (.D(_0030_),
    .CLK(clknet_leaf_35_wb_clk_i),
    .Q(\as2650.stack[3][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8920_ (.D(_0031_),
    .CLK(clknet_leaf_35_wb_clk_i),
    .Q(\as2650.stack[3][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8921_ (.D(_0032_),
    .CLK(clknet_leaf_35_wb_clk_i),
    .Q(\as2650.stack[3][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8922_ (.D(_0033_),
    .CLK(clknet_leaf_54_wb_clk_i),
    .Q(\as2650.stack[3][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8923_ (.D(_0034_),
    .CLK(clknet_leaf_32_wb_clk_i),
    .Q(\as2650.stack[3][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8924_ (.D(_0035_),
    .CLK(clknet_leaf_32_wb_clk_i),
    .Q(\as2650.stack[3][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8925_ (.D(_0036_),
    .CLK(clknet_leaf_32_wb_clk_i),
    .Q(\as2650.stack[3][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8926_ (.D(_0037_),
    .CLK(clknet_leaf_32_wb_clk_i),
    .Q(\as2650.stack[3][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8927_ (.D(_0038_),
    .CLK(clknet_leaf_36_wb_clk_i),
    .Q(\as2650.stack[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8928_ (.D(_0039_),
    .CLK(clknet_leaf_41_wb_clk_i),
    .Q(\as2650.stack[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8929_ (.D(_0040_),
    .CLK(clknet_leaf_41_wb_clk_i),
    .Q(\as2650.stack[2][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8930_ (.D(_0041_),
    .CLK(clknet_leaf_36_wb_clk_i),
    .Q(\as2650.stack[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8931_ (.D(_0042_),
    .CLK(clknet_leaf_32_wb_clk_i),
    .Q(\as2650.stack[2][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8932_ (.D(_0043_),
    .CLK(clknet_leaf_31_wb_clk_i),
    .Q(\as2650.stack[2][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8933_ (.D(_0044_),
    .CLK(clknet_leaf_31_wb_clk_i),
    .Q(\as2650.stack[2][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8934_ (.D(_0045_),
    .CLK(clknet_leaf_31_wb_clk_i),
    .Q(\as2650.stack[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8935_ (.D(_0046_),
    .CLK(clknet_leaf_57_wb_clk_i),
    .Q(\as2650.stack[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8936_ (.D(_0047_),
    .CLK(clknet_leaf_55_wb_clk_i),
    .Q(\as2650.stack[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8937_ (.D(_0048_),
    .CLK(clknet_leaf_55_wb_clk_i),
    .Q(\as2650.stack[1][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8938_ (.D(_0049_),
    .CLK(clknet_leaf_55_wb_clk_i),
    .Q(\as2650.stack[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8939_ (.D(_0050_),
    .CLK(clknet_leaf_58_wb_clk_i),
    .Q(\as2650.stack[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8940_ (.D(_0051_),
    .CLK(clknet_leaf_58_wb_clk_i),
    .Q(\as2650.stack[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8941_ (.D(_0052_),
    .CLK(clknet_leaf_58_wb_clk_i),
    .Q(\as2650.stack[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8942_ (.D(_0053_),
    .CLK(clknet_leaf_58_wb_clk_i),
    .Q(\as2650.stack[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8943_ (.D(_0054_),
    .CLK(clknet_leaf_50_wb_clk_i),
    .Q(\as2650.stack[1][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8944_ (.D(_0055_),
    .CLK(clknet_leaf_51_wb_clk_i),
    .Q(\as2650.stack[1][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8945_ (.D(_0056_),
    .CLK(clknet_leaf_59_wb_clk_i),
    .Q(\as2650.stack[1][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8946_ (.D(_0057_),
    .CLK(clknet_leaf_59_wb_clk_i),
    .Q(\as2650.stack[1][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8947_ (.D(_0058_),
    .CLK(clknet_leaf_50_wb_clk_i),
    .Q(\as2650.stack[1][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8948_ (.D(_0059_),
    .CLK(clknet_leaf_48_wb_clk_i),
    .Q(\as2650.stack[1][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8949_ (.D(_0060_),
    .CLK(clknet_leaf_48_wb_clk_i),
    .Q(\as2650.stack[1][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8950_ (.D(_0061_),
    .CLK(clknet_leaf_54_wb_clk_i),
    .Q(\as2650.stack[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8951_ (.D(_0062_),
    .CLK(clknet_leaf_54_wb_clk_i),
    .Q(\as2650.stack[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8952_ (.D(_0063_),
    .CLK(clknet_leaf_54_wb_clk_i),
    .Q(\as2650.stack[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8953_ (.D(_0064_),
    .CLK(clknet_leaf_54_wb_clk_i),
    .Q(\as2650.stack[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8954_ (.D(_0065_),
    .CLK(clknet_leaf_33_wb_clk_i),
    .Q(\as2650.stack[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8955_ (.D(_0066_),
    .CLK(clknet_leaf_57_wb_clk_i),
    .Q(\as2650.stack[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8956_ (.D(_0067_),
    .CLK(clknet_leaf_57_wb_clk_i),
    .Q(\as2650.stack[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8957_ (.D(_0068_),
    .CLK(clknet_leaf_57_wb_clk_i),
    .Q(\as2650.stack[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8958_ (.D(_0069_),
    .CLK(clknet_leaf_61_wb_clk_i),
    .Q(\as2650.r123_2[3][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8959_ (.D(_0070_),
    .CLK(clknet_leaf_66_wb_clk_i),
    .Q(\as2650.r123_2[3][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8960_ (.D(_0071_),
    .CLK(clknet_leaf_75_wb_clk_i),
    .Q(\as2650.r123_2[3][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8961_ (.D(_0072_),
    .CLK(clknet_3_5__leaf_wb_clk_i),
    .Q(\as2650.r123_2[3][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8962_ (.D(_0073_),
    .CLK(clknet_3_5__leaf_wb_clk_i),
    .Q(\as2650.r123_2[3][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8963_ (.D(_0074_),
    .CLK(clknet_3_5__leaf_wb_clk_i),
    .Q(\as2650.r123_2[3][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8964_ (.D(_0075_),
    .CLK(clknet_leaf_61_wb_clk_i),
    .Q(\as2650.r123_2[3][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8965_ (.D(_0076_),
    .CLK(clknet_leaf_63_wb_clk_i),
    .Q(\as2650.r123_2[3][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8966_ (.D(_0077_),
    .CLK(clknet_leaf_43_wb_clk_i),
    .Q(\as2650.psu[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8967_ (.D(_0078_),
    .CLK(clknet_leaf_15_wb_clk_i),
    .Q(net42));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8968_ (.D(_0079_),
    .CLK(clknet_leaf_15_wb_clk_i),
    .Q(net43));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8969_ (.D(_0080_),
    .CLK(clknet_leaf_15_wb_clk_i),
    .Q(net44));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8970_ (.D(_0081_),
    .CLK(clknet_leaf_15_wb_clk_i),
    .Q(net45));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8971_ (.D(_0082_),
    .CLK(clknet_leaf_15_wb_clk_i),
    .Q(net46));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8972_ (.D(_0083_),
    .CLK(clknet_leaf_15_wb_clk_i),
    .Q(net20));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8973_ (.D(_0084_),
    .CLK(clknet_leaf_16_wb_clk_i),
    .Q(net21));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8974_ (.D(_0085_),
    .CLK(clknet_leaf_16_wb_clk_i),
    .Q(net22));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8975_ (.D(_0086_),
    .CLK(clknet_leaf_47_wb_clk_i),
    .Q(\as2650.stack[3][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8976_ (.D(_0087_),
    .CLK(clknet_leaf_51_wb_clk_i),
    .Q(\as2650.stack[3][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8977_ (.D(_0088_),
    .CLK(clknet_leaf_51_wb_clk_i),
    .Q(\as2650.stack[3][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8978_ (.D(_0089_),
    .CLK(clknet_leaf_51_wb_clk_i),
    .Q(\as2650.stack[3][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8979_ (.D(_0090_),
    .CLK(clknet_leaf_50_wb_clk_i),
    .Q(\as2650.stack[3][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8980_ (.D(_0091_),
    .CLK(clknet_leaf_48_wb_clk_i),
    .Q(\as2650.stack[3][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8981_ (.D(_0092_),
    .CLK(clknet_leaf_47_wb_clk_i),
    .Q(\as2650.stack[3][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8982_ (.D(_0093_),
    .CLK(clknet_3_1__leaf_wb_clk_i),
    .Q(\as2650.psl[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8983_ (.D(_0094_),
    .CLK(clknet_leaf_69_wb_clk_i),
    .Q(\as2650.psl[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8984_ (.D(_0095_),
    .CLK(clknet_leaf_7_wb_clk_i),
    .Q(\as2650.ins_reg[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8985_ (.D(_0096_),
    .CLK(clknet_leaf_7_wb_clk_i),
    .Q(\as2650.ins_reg[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8986_ (.D(_0097_),
    .CLK(clknet_leaf_3_wb_clk_i),
    .Q(\as2650.ins_reg[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8987_ (.D(_0098_),
    .CLK(clknet_leaf_1_wb_clk_i),
    .Q(\as2650.alu_op[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8988_ (.D(_0099_),
    .CLK(clknet_leaf_9_wb_clk_i),
    .Q(\as2650.alu_op[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8989_ (.D(_0100_),
    .CLK(clknet_leaf_9_wb_clk_i),
    .Q(\as2650.alu_op[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8990_ (.D(_0101_),
    .CLK(clknet_leaf_50_wb_clk_i),
    .Q(\as2650.stack[0][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8991_ (.D(_0102_),
    .CLK(clknet_leaf_51_wb_clk_i),
    .Q(\as2650.stack[0][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8992_ (.D(_0103_),
    .CLK(clknet_leaf_59_wb_clk_i),
    .Q(\as2650.stack[0][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8993_ (.D(_0104_),
    .CLK(clknet_leaf_59_wb_clk_i),
    .Q(\as2650.stack[0][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8994_ (.D(_0105_),
    .CLK(clknet_leaf_50_wb_clk_i),
    .Q(\as2650.stack[0][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8995_ (.D(_0106_),
    .CLK(clknet_leaf_67_wb_clk_i),
    .Q(\as2650.stack[0][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8996_ (.D(_0107_),
    .CLK(clknet_leaf_49_wb_clk_i),
    .Q(\as2650.stack[0][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8997_ (.D(_0108_),
    .CLK(clknet_leaf_47_wb_clk_i),
    .Q(\as2650.stack[6][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8998_ (.D(_0109_),
    .CLK(clknet_leaf_52_wb_clk_i),
    .Q(\as2650.stack[6][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8999_ (.D(_0110_),
    .CLK(clknet_leaf_52_wb_clk_i),
    .Q(\as2650.stack[6][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9000_ (.D(_0111_),
    .CLK(clknet_leaf_53_wb_clk_i),
    .Q(\as2650.stack[6][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9001_ (.D(_0112_),
    .CLK(clknet_leaf_46_wb_clk_i),
    .Q(\as2650.stack[6][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9002_ (.D(_0113_),
    .CLK(clknet_leaf_48_wb_clk_i),
    .Q(\as2650.stack[6][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9003_ (.D(_0114_),
    .CLK(clknet_leaf_44_wb_clk_i),
    .Q(\as2650.stack[6][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9004_ (.D(_0115_),
    .CLK(clknet_leaf_77_wb_clk_i),
    .Q(\as2650.r123_2[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9005_ (.D(_0116_),
    .CLK(clknet_leaf_79_wb_clk_i),
    .Q(\as2650.r123_2[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9006_ (.D(_0117_),
    .CLK(clknet_leaf_78_wb_clk_i),
    .Q(\as2650.r123_2[2][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9007_ (.D(_0118_),
    .CLK(clknet_leaf_78_wb_clk_i),
    .Q(\as2650.r123_2[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9008_ (.D(_0119_),
    .CLK(clknet_leaf_1_wb_clk_i),
    .Q(\as2650.r123_2[2][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9009_ (.D(_0120_),
    .CLK(clknet_leaf_78_wb_clk_i),
    .Q(\as2650.r123_2[2][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9010_ (.D(_0121_),
    .CLK(clknet_leaf_77_wb_clk_i),
    .Q(\as2650.r123_2[2][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9011_ (.D(_0122_),
    .CLK(clknet_leaf_77_wb_clk_i),
    .Q(\as2650.r123_2[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9012_ (.D(_0123_),
    .CLK(clknet_leaf_34_wb_clk_i),
    .Q(\as2650.stack[5][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9013_ (.D(_0124_),
    .CLK(clknet_leaf_35_wb_clk_i),
    .Q(\as2650.stack[5][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9014_ (.D(_0125_),
    .CLK(clknet_leaf_34_wb_clk_i),
    .Q(\as2650.stack[5][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9015_ (.D(_0126_),
    .CLK(clknet_leaf_35_wb_clk_i),
    .Q(\as2650.stack[5][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9016_ (.D(_0127_),
    .CLK(clknet_leaf_30_wb_clk_i),
    .Q(\as2650.stack[5][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9017_ (.D(_0128_),
    .CLK(clknet_leaf_30_wb_clk_i),
    .Q(\as2650.stack[5][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9018_ (.D(_0129_),
    .CLK(clknet_leaf_31_wb_clk_i),
    .Q(\as2650.stack[5][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9019_ (.D(_0130_),
    .CLK(clknet_leaf_31_wb_clk_i),
    .Q(\as2650.stack[5][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9020_ (.D(_0131_),
    .CLK(clknet_leaf_74_wb_clk_i),
    .Q(\as2650.r123_2[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9021_ (.D(_0132_),
    .CLK(clknet_leaf_5_wb_clk_i),
    .Q(\as2650.r123_2[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9022_ (.D(_0133_),
    .CLK(clknet_leaf_5_wb_clk_i),
    .Q(\as2650.r123_2[1][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9023_ (.D(_0134_),
    .CLK(clknet_leaf_74_wb_clk_i),
    .Q(\as2650.r123_2[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9024_ (.D(_0135_),
    .CLK(clknet_leaf_5_wb_clk_i),
    .Q(\as2650.r123_2[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9025_ (.D(_0136_),
    .CLK(clknet_leaf_71_wb_clk_i),
    .Q(\as2650.r123_2[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9026_ (.D(_0137_),
    .CLK(clknet_leaf_74_wb_clk_i),
    .Q(\as2650.r123_2[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9027_ (.D(_0138_),
    .CLK(clknet_leaf_73_wb_clk_i),
    .Q(\as2650.r123_2[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9028_ (.D(_0139_),
    .CLK(clknet_leaf_20_wb_clk_i),
    .Q(\as2650.addr_buff[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9029_ (.D(_0140_),
    .CLK(clknet_leaf_20_wb_clk_i),
    .Q(\as2650.addr_buff[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9030_ (.D(_0141_),
    .CLK(clknet_leaf_20_wb_clk_i),
    .Q(\as2650.addr_buff[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9031_ (.D(_0142_),
    .CLK(clknet_leaf_20_wb_clk_i),
    .Q(\as2650.addr_buff[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9032_ (.D(_0143_),
    .CLK(clknet_leaf_21_wb_clk_i),
    .Q(\as2650.addr_buff[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9033_ (.D(_0144_),
    .CLK(clknet_leaf_9_wb_clk_i),
    .Q(\as2650.addr_buff[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9034_ (.D(_0145_),
    .CLK(clknet_leaf_9_wb_clk_i),
    .Q(\as2650.addr_buff[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9035_ (.D(_0146_),
    .CLK(clknet_leaf_13_wb_clk_i),
    .Q(\as2650.addr_buff[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9036_ (.D(_0000_),
    .CLK(clknet_leaf_18_wb_clk_i),
    .Q(\as2650.cycle[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9037_ (.D(_0005_),
    .CLK(clknet_leaf_13_wb_clk_i),
    .Q(\as2650.cycle[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9038_ (.D(_0006_),
    .CLK(clknet_leaf_14_wb_clk_i),
    .Q(\as2650.cycle[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9039_ (.D(_0007_),
    .CLK(clknet_leaf_13_wb_clk_i),
    .Q(\as2650.cycle[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9040_ (.D(_0008_),
    .CLK(clknet_3_2__leaf_wb_clk_i),
    .Q(\as2650.cycle[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9041_ (.D(_0009_),
    .CLK(clknet_leaf_13_wb_clk_i),
    .Q(\as2650.cycle[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9042_ (.D(_0010_),
    .CLK(clknet_leaf_40_wb_clk_i),
    .Q(\as2650.cycle[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9043_ (.D(_0011_),
    .CLK(clknet_leaf_15_wb_clk_i),
    .Q(\as2650.cycle[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9044_ (.D(_0012_),
    .CLK(clknet_leaf_21_wb_clk_i),
    .Q(\as2650.cycle[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9045_ (.D(_0013_),
    .CLK(clknet_leaf_13_wb_clk_i),
    .Q(\as2650.cycle[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9046_ (.D(_0001_),
    .CLK(clknet_leaf_14_wb_clk_i),
    .Q(\as2650.cycle[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9047_ (.D(_0002_),
    .CLK(clknet_3_2__leaf_wb_clk_i),
    .Q(\as2650.cycle[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9048_ (.D(_0003_),
    .CLK(clknet_leaf_14_wb_clk_i),
    .Q(\as2650.cycle[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9049_ (.D(_0004_),
    .CLK(clknet_leaf_29_wb_clk_i),
    .Q(\as2650.cycle[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9050_ (.D(_0147_),
    .CLK(clknet_leaf_46_wb_clk_i),
    .Q(\as2650.stack[4][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9051_ (.D(_0148_),
    .CLK(clknet_leaf_54_wb_clk_i),
    .Q(\as2650.stack[4][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9052_ (.D(_0149_),
    .CLK(clknet_leaf_56_wb_clk_i),
    .Q(\as2650.stack[4][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9053_ (.D(_0150_),
    .CLK(clknet_leaf_53_wb_clk_i),
    .Q(\as2650.stack[4][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9054_ (.D(_0151_),
    .CLK(clknet_leaf_46_wb_clk_i),
    .Q(\as2650.stack[4][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9055_ (.D(_0152_),
    .CLK(clknet_leaf_45_wb_clk_i),
    .Q(\as2650.stack[4][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9056_ (.D(_0153_),
    .CLK(clknet_leaf_44_wb_clk_i),
    .Q(\as2650.stack[4][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9057_ (.D(_0154_),
    .CLK(clknet_leaf_70_wb_clk_i),
    .Q(\as2650.r123_2[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9058_ (.D(_0155_),
    .CLK(clknet_leaf_70_wb_clk_i),
    .Q(\as2650.r123_2[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9059_ (.D(_0156_),
    .CLK(clknet_leaf_70_wb_clk_i),
    .Q(\as2650.r123_2[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9060_ (.D(_0157_),
    .CLK(clknet_leaf_70_wb_clk_i),
    .Q(\as2650.r123_2[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9061_ (.D(_0158_),
    .CLK(clknet_leaf_70_wb_clk_i),
    .Q(\as2650.r123_2[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9062_ (.D(_0159_),
    .CLK(clknet_leaf_70_wb_clk_i),
    .Q(\as2650.r123_2[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9063_ (.D(_0160_),
    .CLK(clknet_leaf_70_wb_clk_i),
    .Q(\as2650.r123_2[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9064_ (.D(_0161_),
    .CLK(clknet_leaf_70_wb_clk_i),
    .Q(\as2650.r123_2[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9065_ (.D(_0162_),
    .CLK(clknet_leaf_49_wb_clk_i),
    .Q(\as2650.stack[2][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9066_ (.D(_0163_),
    .CLK(clknet_leaf_51_wb_clk_i),
    .Q(\as2650.stack[2][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9067_ (.D(_0164_),
    .CLK(clknet_leaf_52_wb_clk_i),
    .Q(\as2650.stack[2][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9068_ (.D(_0165_),
    .CLK(clknet_leaf_59_wb_clk_i),
    .Q(\as2650.stack[2][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9069_ (.D(_0166_),
    .CLK(clknet_leaf_50_wb_clk_i),
    .Q(\as2650.stack[2][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9070_ (.D(_0167_),
    .CLK(clknet_leaf_48_wb_clk_i),
    .Q(\as2650.stack[2][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9071_ (.D(_0168_),
    .CLK(clknet_leaf_48_wb_clk_i),
    .Q(\as2650.stack[2][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9072_ (.D(_0169_),
    .CLK(clknet_leaf_17_wb_clk_i),
    .Q(net25));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9073_ (.D(_0170_),
    .CLK(clknet_leaf_17_wb_clk_i),
    .Q(net23));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9074_ (.D(_0171_),
    .CLK(clknet_leaf_18_wb_clk_i),
    .Q(net24));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9075_ (.D(_0172_),
    .CLK(clknet_leaf_19_wb_clk_i),
    .Q(net29));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9076_ (.D(_0173_),
    .CLK(clknet_leaf_19_wb_clk_i),
    .Q(net30));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9077_ (.D(_0174_),
    .CLK(clknet_leaf_19_wb_clk_i),
    .Q(net31));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9078_ (.D(_0175_),
    .CLK(clknet_leaf_22_wb_clk_i),
    .Q(net32));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9079_ (.D(_0176_),
    .CLK(clknet_leaf_19_wb_clk_i),
    .Q(net33));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9080_ (.D(_0177_),
    .CLK(clknet_leaf_23_wb_clk_i),
    .Q(net34));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9081_ (.D(_0178_),
    .CLK(clknet_leaf_22_wb_clk_i),
    .Q(net35));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9082_ (.D(_0179_),
    .CLK(clknet_leaf_22_wb_clk_i),
    .Q(net36));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9083_ (.D(_0180_),
    .CLK(clknet_leaf_22_wb_clk_i),
    .Q(net37));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9084_ (.D(_0181_),
    .CLK(clknet_leaf_23_wb_clk_i),
    .Q(net38));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9085_ (.D(_0182_),
    .CLK(clknet_leaf_23_wb_clk_i),
    .Q(net39));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9086_ (.D(_0183_),
    .CLK(clknet_leaf_23_wb_clk_i),
    .Q(net40));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9087_ (.D(_0184_),
    .CLK(clknet_leaf_23_wb_clk_i),
    .Q(net41));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9088_ (.D(_0185_),
    .CLK(clknet_leaf_16_wb_clk_i),
    .Q(net27));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9089_ (.D(_0186_),
    .CLK(clknet_leaf_17_wb_clk_i),
    .Q(net26));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9090_ (.D(_0187_),
    .CLK(clknet_leaf_9_wb_clk_i),
    .Q(\as2650.idx_ctrl[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9091_ (.D(_0188_),
    .CLK(clknet_leaf_9_wb_clk_i),
    .Q(\as2650.idx_ctrl[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9092_ (.D(_0189_),
    .CLK(clknet_leaf_81_wb_clk_i),
    .Q(\as2650.holding_reg[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9093_ (.D(_0190_),
    .CLK(clknet_leaf_1_wb_clk_i),
    .Q(\as2650.holding_reg[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9094_ (.D(_0191_),
    .CLK(clknet_leaf_82_wb_clk_i),
    .Q(\as2650.holding_reg[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9095_ (.D(_0192_),
    .CLK(clknet_3_0__leaf_wb_clk_i),
    .Q(\as2650.holding_reg[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9096_ (.D(_0193_),
    .CLK(clknet_leaf_1_wb_clk_i),
    .Q(\as2650.holding_reg[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9097_ (.D(_0194_),
    .CLK(clknet_leaf_82_wb_clk_i),
    .Q(\as2650.holding_reg[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9098_ (.D(_0195_),
    .CLK(clknet_leaf_82_wb_clk_i),
    .Q(\as2650.holding_reg[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9099_ (.D(_0196_),
    .CLK(clknet_leaf_82_wb_clk_i),
    .Q(\as2650.holding_reg[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9100_ (.D(_0197_),
    .CLK(clknet_leaf_37_wb_clk_i),
    .Q(\as2650.halted ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9101_ (.D(_0198_),
    .CLK(clknet_leaf_40_wb_clk_i),
    .Q(\as2650.psu[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9102_ (.D(_0199_),
    .CLK(clknet_leaf_15_wb_clk_i),
    .Q(\as2650.pc[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9103_ (.D(_0200_),
    .CLK(clknet_3_6__leaf_wb_clk_i),
    .Q(\as2650.pc[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9104_ (.D(_0201_),
    .CLK(clknet_leaf_27_wb_clk_i),
    .Q(\as2650.pc[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9105_ (.D(_0202_),
    .CLK(clknet_leaf_25_wb_clk_i),
    .Q(\as2650.pc[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9106_ (.D(_0203_),
    .CLK(clknet_leaf_25_wb_clk_i),
    .Q(\as2650.pc[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9107_ (.D(_0204_),
    .CLK(clknet_leaf_24_wb_clk_i),
    .Q(\as2650.pc[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9108_ (.D(_0205_),
    .CLK(clknet_leaf_25_wb_clk_i),
    .Q(\as2650.pc[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9109_ (.D(_0206_),
    .CLK(clknet_leaf_27_wb_clk_i),
    .Q(\as2650.pc[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9110_ (.D(_0207_),
    .CLK(clknet_leaf_24_wb_clk_i),
    .Q(\as2650.pc[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9111_ (.D(_0208_),
    .CLK(clknet_leaf_27_wb_clk_i),
    .Q(\as2650.pc[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9112_ (.D(_0209_),
    .CLK(clknet_leaf_27_wb_clk_i),
    .Q(\as2650.pc[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9113_ (.D(_0210_),
    .CLK(clknet_3_6__leaf_wb_clk_i),
    .Q(\as2650.pc[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9114_ (.D(_0211_),
    .CLK(clknet_leaf_29_wb_clk_i),
    .Q(\as2650.pc[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9115_ (.D(_0212_),
    .CLK(clknet_leaf_38_wb_clk_i),
    .Q(\as2650.pc[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9116_ (.D(_0213_),
    .CLK(clknet_3_6__leaf_wb_clk_i),
    .Q(\as2650.pc[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9117_ (.D(_0214_),
    .CLK(clknet_leaf_80_wb_clk_i),
    .Q(\as2650.r0[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9118_ (.D(_0215_),
    .CLK(clknet_leaf_80_wb_clk_i),
    .Q(\as2650.r0[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9119_ (.D(_0216_),
    .CLK(clknet_leaf_80_wb_clk_i),
    .Q(\as2650.r0[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9120_ (.D(_0217_),
    .CLK(clknet_leaf_80_wb_clk_i),
    .Q(\as2650.r0[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9121_ (.D(_0218_),
    .CLK(clknet_leaf_81_wb_clk_i),
    .Q(\as2650.r0[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9122_ (.D(_0219_),
    .CLK(clknet_leaf_81_wb_clk_i),
    .Q(\as2650.r0[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9123_ (.D(_0220_),
    .CLK(clknet_leaf_82_wb_clk_i),
    .Q(\as2650.r0[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9124_ (.D(_0221_),
    .CLK(clknet_leaf_81_wb_clk_i),
    .Q(\as2650.r0[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9125_ (.D(_0222_),
    .CLK(clknet_leaf_34_wb_clk_i),
    .Q(\as2650.stack[7][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9126_ (.D(_0223_),
    .CLK(clknet_leaf_38_wb_clk_i),
    .Q(\as2650.stack[7][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9127_ (.D(_0224_),
    .CLK(clknet_leaf_38_wb_clk_i),
    .Q(\as2650.stack[7][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9128_ (.D(_0225_),
    .CLK(clknet_leaf_34_wb_clk_i),
    .Q(\as2650.stack[7][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9129_ (.D(_0226_),
    .CLK(clknet_leaf_33_wb_clk_i),
    .Q(\as2650.stack[7][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9130_ (.D(_0227_),
    .CLK(clknet_leaf_33_wb_clk_i),
    .Q(\as2650.stack[7][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9131_ (.D(_0228_),
    .CLK(clknet_leaf_30_wb_clk_i),
    .Q(\as2650.stack[7][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9132_ (.D(_0229_),
    .CLK(clknet_leaf_33_wb_clk_i),
    .Q(\as2650.stack[7][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9133_ (.D(_0230_),
    .CLK(clknet_leaf_46_wb_clk_i),
    .Q(\as2650.stack[7][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9134_ (.D(_0231_),
    .CLK(clknet_leaf_56_wb_clk_i),
    .Q(\as2650.stack[7][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9135_ (.D(_0232_),
    .CLK(clknet_leaf_56_wb_clk_i),
    .Q(\as2650.stack[7][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9136_ (.D(_0233_),
    .CLK(clknet_leaf_53_wb_clk_i),
    .Q(\as2650.stack[7][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9137_ (.D(_0234_),
    .CLK(clknet_leaf_53_wb_clk_i),
    .Q(\as2650.stack[7][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9138_ (.D(_0235_),
    .CLK(clknet_leaf_44_wb_clk_i),
    .Q(\as2650.stack[7][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9139_ (.D(_0236_),
    .CLK(clknet_leaf_44_wb_clk_i),
    .Q(\as2650.stack[7][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9140_ (.D(_0237_),
    .CLK(clknet_leaf_37_wb_clk_i),
    .Q(\as2650.stack[6][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9141_ (.D(_0238_),
    .CLK(clknet_leaf_37_wb_clk_i),
    .Q(\as2650.stack[6][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9142_ (.D(_0239_),
    .CLK(clknet_leaf_37_wb_clk_i),
    .Q(\as2650.stack[6][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9143_ (.D(_0240_),
    .CLK(clknet_leaf_37_wb_clk_i),
    .Q(\as2650.stack[6][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9144_ (.D(_0241_),
    .CLK(clknet_leaf_30_wb_clk_i),
    .Q(\as2650.stack[6][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9145_ (.D(_0242_),
    .CLK(clknet_leaf_30_wb_clk_i),
    .Q(\as2650.stack[6][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9146_ (.D(_0243_),
    .CLK(clknet_leaf_34_wb_clk_i),
    .Q(\as2650.stack[6][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9147_ (.D(_0244_),
    .CLK(clknet_leaf_34_wb_clk_i),
    .Q(\as2650.stack[6][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9148_ (.D(_0245_),
    .CLK(clknet_leaf_46_wb_clk_i),
    .Q(\as2650.stack[5][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9149_ (.D(_0246_),
    .CLK(clknet_leaf_56_wb_clk_i),
    .Q(\as2650.stack[5][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9150_ (.D(_0247_),
    .CLK(clknet_leaf_56_wb_clk_i),
    .Q(\as2650.stack[5][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9151_ (.D(_0248_),
    .CLK(clknet_leaf_53_wb_clk_i),
    .Q(\as2650.stack[5][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9152_ (.D(_0249_),
    .CLK(clknet_leaf_46_wb_clk_i),
    .Q(\as2650.stack[5][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9153_ (.D(_0250_),
    .CLK(clknet_leaf_45_wb_clk_i),
    .Q(\as2650.stack[5][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9154_ (.D(_0251_),
    .CLK(clknet_leaf_44_wb_clk_i),
    .Q(\as2650.stack[5][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9155_ (.D(_0252_),
    .CLK(clknet_leaf_71_wb_clk_i),
    .Q(\as2650.r123[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9156_ (.D(_0253_),
    .CLK(clknet_leaf_6_wb_clk_i),
    .Q(\as2650.r123[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9157_ (.D(_0254_),
    .CLK(clknet_leaf_3_wb_clk_i),
    .Q(\as2650.r123[1][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9158_ (.D(_0255_),
    .CLK(clknet_leaf_73_wb_clk_i),
    .Q(\as2650.r123[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9159_ (.D(_0256_),
    .CLK(clknet_leaf_6_wb_clk_i),
    .Q(\as2650.r123[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9160_ (.D(_0257_),
    .CLK(clknet_leaf_71_wb_clk_i),
    .Q(\as2650.r123[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9161_ (.D(_0258_),
    .CLK(clknet_leaf_73_wb_clk_i),
    .Q(\as2650.r123[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9162_ (.D(_0259_),
    .CLK(clknet_leaf_71_wb_clk_i),
    .Q(\as2650.r123[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9163_ (.D(_0260_),
    .CLK(clknet_leaf_77_wb_clk_i),
    .Q(\as2650.r123[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9164_ (.D(_0261_),
    .CLK(clknet_leaf_79_wb_clk_i),
    .Q(\as2650.r123[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9165_ (.D(_0262_),
    .CLK(clknet_leaf_2_wb_clk_i),
    .Q(\as2650.r123[2][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9166_ (.D(_0263_),
    .CLK(clknet_leaf_4_wb_clk_i),
    .Q(\as2650.r123[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9167_ (.D(_0264_),
    .CLK(clknet_leaf_2_wb_clk_i),
    .Q(\as2650.r123[2][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9168_ (.D(_0265_),
    .CLK(clknet_leaf_78_wb_clk_i),
    .Q(\as2650.r123[2][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9169_ (.D(_0266_),
    .CLK(clknet_leaf_4_wb_clk_i),
    .Q(\as2650.r123[2][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9170_ (.D(_0267_),
    .CLK(clknet_leaf_5_wb_clk_i),
    .Q(\as2650.r123[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9171_ (.D(_0268_),
    .CLK(clknet_leaf_36_wb_clk_i),
    .Q(\as2650.stack[4][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9172_ (.D(_0269_),
    .CLK(clknet_leaf_36_wb_clk_i),
    .Q(\as2650.stack[4][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9173_ (.D(_0270_),
    .CLK(clknet_leaf_36_wb_clk_i),
    .Q(\as2650.stack[4][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9174_ (.D(_0271_),
    .CLK(clknet_leaf_36_wb_clk_i),
    .Q(\as2650.stack[4][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9175_ (.D(_0272_),
    .CLK(clknet_leaf_31_wb_clk_i),
    .Q(\as2650.stack[4][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9176_ (.D(_0273_),
    .CLK(clknet_leaf_31_wb_clk_i),
    .Q(\as2650.stack[4][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9177_ (.D(_0274_),
    .CLK(clknet_leaf_31_wb_clk_i),
    .Q(\as2650.stack[4][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9178_ (.D(_0275_),
    .CLK(clknet_leaf_31_wb_clk_i),
    .Q(\as2650.stack[4][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9179_ (.D(_0276_),
    .CLK(clknet_leaf_69_wb_clk_i),
    .Q(\as2650.ins_reg[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9180_ (.D(_0277_),
    .CLK(clknet_3_2__leaf_wb_clk_i),
    .Q(\as2650.ins_reg[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9181_ (.D(_0278_),
    .CLK(clknet_leaf_45_wb_clk_i),
    .Q(\as2650.psu[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9182_ (.D(_0279_),
    .CLK(clknet_leaf_41_wb_clk_i),
    .Q(\as2650.psu[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9183_ (.D(_0280_),
    .CLK(clknet_leaf_41_wb_clk_i),
    .Q(\as2650.psu[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9184_ (.D(_0281_),
    .CLK(clknet_leaf_82_wb_clk_i),
    .Q(\as2650.carry ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9185_ (.D(_0282_),
    .CLK(clknet_3_7__leaf_wb_clk_i),
    .Q(\as2650.psl[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9186_ (.D(_0283_),
    .CLK(clknet_leaf_44_wb_clk_i),
    .Q(\as2650.overflow ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9187_ (.D(_0284_),
    .CLK(clknet_leaf_67_wb_clk_i),
    .Q(\as2650.psl[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9188_ (.D(_0285_),
    .CLK(clknet_leaf_44_wb_clk_i),
    .Q(\as2650.psl[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9189_ (.D(_0286_),
    .CLK(clknet_leaf_43_wb_clk_i),
    .Q(\as2650.psl[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9190_ (.D(_0287_),
    .CLK(clknet_leaf_43_wb_clk_i),
    .Q(net28));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9191_ (.D(_0288_),
    .CLK(clknet_leaf_45_wb_clk_i),
    .Q(\as2650.psu[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9192_ (.D(_0289_),
    .CLK(clknet_leaf_45_wb_clk_i),
    .Q(\as2650.psu[3] ));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_87 (.Z(net87));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_88 (.Z(net88));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_89 (.Z(net89));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_90 (.Z(net90));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_91 (.Z(net91));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_92 (.Z(net92));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_93 (.Z(net93));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_94 (.Z(net94));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_95 (.Z(net95));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_96 (.Z(net96));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_1_wb_clk_i (.I(clknet_3_2__leaf_wb_clk_i),
    .Z(clknet_leaf_1_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_57 (.ZN(net57));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_58 (.ZN(net58));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_59 (.ZN(net59));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_60 (.ZN(net60));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_61 (.ZN(net61));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_62 (.ZN(net62));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_63 (.ZN(net63));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_64 (.ZN(net64));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_65 (.ZN(net65));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_66 (.ZN(net66));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_67 (.ZN(net67));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_68 (.ZN(net68));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_69 (.ZN(net69));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_70 (.ZN(net70));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_71 (.ZN(net71));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_72 (.ZN(net72));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_73 (.ZN(net73));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_74 (.ZN(net74));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_75 (.ZN(net75));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_76 (.ZN(net76));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_77 (.ZN(net77));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_78 (.ZN(net78));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_79 (.ZN(net79));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_80 (.ZN(net80));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_81 (.ZN(net81));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_82 (.ZN(net82));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_83 (.ZN(net83));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_84 (.ZN(net84));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_85 (.ZN(net85));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_86 (.Z(net86));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _9234_ (.I(net47),
    .Z(net15));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _9235_ (.I(net47),
    .Z(net16));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _9236_ (.I(net47),
    .Z(net17));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _9237_ (.I(net47),
    .Z(net18));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _9238_ (.I(net48),
    .Z(net19));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _9239_ (.I(net48),
    .Z(net12));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _9240_ (.I(net48),
    .Z(net13));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_0 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_7 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_8 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_9 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_10 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_11 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_12 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_13 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_14 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_15 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_16 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_17 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_18 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_19 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_20 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_21 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_22 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_23 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_24 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_25 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_26 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_27 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_28 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_29 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_30 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_31 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_32 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_33 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_34 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_35 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_36 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_37 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_38 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_39 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_40 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_41 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_42 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_43 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_44 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_45 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_46 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_47 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_48 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_49 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_50 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_51 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_52 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_53 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_54 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_55 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_56 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_57 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_58 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_59 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_60 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_61 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_62 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_63 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_64 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_65 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_66 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_67 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_68 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_69 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_70 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_71 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_72 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_73 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_74 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_75 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_76 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_77 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_78 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_79 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_80 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_81 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_82 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_83 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_84 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_85 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_86 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_87 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_88 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_89 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_90 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_91 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_92 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_93 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_94 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_95 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_96 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_97 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_98 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_99 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_100 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_101 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_102 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_103 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_104 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_105 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_106 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_107 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_108 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_109 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_110 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_111 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_112 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_113 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_114 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_115 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_116 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_117 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_118 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_119 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_120 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_121 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_122 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_123 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_124 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_125 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_126 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_127 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_128 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_129 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_130 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_131 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_132 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_133 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_134 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_135 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_136 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_137 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_138 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_139 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_140 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_141 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_142 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_143 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_144 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_145 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_146 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_147 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_148 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_149 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_150 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_151 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_152 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_153 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_154 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_155 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_156 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_157 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_158 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_159 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_160 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_161 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_162 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_163 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_164 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_165 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_166 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_167 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_168 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_169 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_170 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_171 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_172 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_173 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_174 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_175 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_176 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_177 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_178 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_179 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_180 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_181 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_182 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_183 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_184 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_185 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_186 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_187 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_188 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_189 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_190 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_191 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_192 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_193 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_194 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_195 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_196 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_197 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_198 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_199 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_200 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_201 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_202 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_203 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_204 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_205 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_206 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_207 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_208 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_209 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_210 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_211 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_212 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_213 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_214 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_215 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_216 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_217 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_218 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_219 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_220 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_221 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_222 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_223 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_224 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_225 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_226 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_227 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_228 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_229 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_230 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_231 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_232 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_233 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_234 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_235 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_236 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_237 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_238 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_239 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_240 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_241 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_242 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_243 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_244 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_245 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_246 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_247 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_248 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_249 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_250 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_251 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_252 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_253 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_254 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_255 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_256 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_257 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_258 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_259 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_260 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_261 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_262 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_263 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_264 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_265 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_266 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_267 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_268 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_269 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_270 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_271 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_272 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_273 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_274 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_275 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_276 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_277 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_278 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_279 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_280 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_281 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_282 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_283 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_284 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_285 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_286 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_287 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_288 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3525 ();
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input1 (.I(io_in[10]),
    .Z(net1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input2 (.I(io_in[11]),
    .Z(net2));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input3 (.I(io_in[12]),
    .Z(net3));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input4 (.I(io_in[13]),
    .Z(net4));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input5 (.I(io_in[33]),
    .Z(net5));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input6 (.I(io_in[34]),
    .Z(net6));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input7 (.I(io_in[5]),
    .Z(net7));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input8 (.I(io_in[6]),
    .Z(net8));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input9 (.I(io_in[7]),
    .Z(net9));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input10 (.I(io_in[8]),
    .Z(net10));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input11 (.I(io_in[9]),
    .Z(net11));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output12 (.I(net12),
    .Z(io_oeb[10]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output13 (.I(net13),
    .Z(io_oeb[11]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output14 (.I(net51),
    .Z(io_oeb[12]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output15 (.I(net15),
    .Z(io_oeb[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output16 (.I(net16),
    .Z(io_oeb[6]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output17 (.I(net17),
    .Z(io_oeb[7]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output18 (.I(net18),
    .Z(io_oeb[8]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output19 (.I(net19),
    .Z(io_oeb[9]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output20 (.I(net20),
    .Z(io_out[10]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output21 (.I(net21),
    .Z(io_out[11]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output22 (.I(net22),
    .Z(io_out[12]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output23 (.I(net23),
    .Z(io_out[14]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output24 (.I(net24),
    .Z(io_out[15]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output25 (.I(net25),
    .Z(io_out[16]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output26 (.I(net26),
    .Z(io_out[17]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output27 (.I(net27),
    .Z(io_out[18]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output28 (.I(net28),
    .Z(io_out[19]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output29 (.I(net29),
    .Z(io_out[20]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output30 (.I(net30),
    .Z(io_out[21]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output31 (.I(net31),
    .Z(io_out[22]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output32 (.I(net32),
    .Z(io_out[23]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output33 (.I(net33),
    .Z(io_out[24]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output34 (.I(net34),
    .Z(io_out[25]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output35 (.I(net35),
    .Z(io_out[26]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output36 (.I(net36),
    .Z(io_out[27]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output37 (.I(net37),
    .Z(io_out[28]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output38 (.I(net38),
    .Z(io_out[29]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output39 (.I(net39),
    .Z(io_out[30]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output40 (.I(net40),
    .Z(io_out[31]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output41 (.I(net41),
    .Z(io_out[32]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output42 (.I(net42),
    .Z(io_out[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output43 (.I(net43),
    .Z(io_out[6]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output44 (.I(net44),
    .Z(io_out[7]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output45 (.I(net45),
    .Z(io_out[8]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output46 (.I(net46),
    .Z(io_out[9]));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout47 (.I(net49),
    .Z(net47));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout48 (.I(net49),
    .Z(net48));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout49 (.I(net50),
    .Z(net49));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout50 (.I(net51),
    .Z(net50));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout51 (.I(net14),
    .Z(net51));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout52 (.I(net26),
    .Z(net52));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout53 (.I(net41),
    .Z(net53));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout54 (.I(net36),
    .Z(net54));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout55 (.I(net32),
    .Z(net55));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_56 (.ZN(net56));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_2_wb_clk_i (.I(clknet_3_0__leaf_wb_clk_i),
    .Z(clknet_leaf_2_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_3_wb_clk_i (.I(clknet_opt_1_0_wb_clk_i),
    .Z(clknet_leaf_3_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_4_wb_clk_i (.I(clknet_3_0__leaf_wb_clk_i),
    .Z(clknet_leaf_4_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_5_wb_clk_i (.I(clknet_3_1__leaf_wb_clk_i),
    .Z(clknet_leaf_5_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_6_wb_clk_i (.I(clknet_3_1__leaf_wb_clk_i),
    .Z(clknet_leaf_6_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_7_wb_clk_i (.I(clknet_3_1__leaf_wb_clk_i),
    .Z(clknet_leaf_7_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_9_wb_clk_i (.I(clknet_3_2__leaf_wb_clk_i),
    .Z(clknet_leaf_9_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_13_wb_clk_i (.I(clknet_3_2__leaf_wb_clk_i),
    .Z(clknet_leaf_13_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_14_wb_clk_i (.I(clknet_3_2__leaf_wb_clk_i),
    .Z(clknet_leaf_14_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_15_wb_clk_i (.I(clknet_3_2__leaf_wb_clk_i),
    .Z(clknet_leaf_15_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_16_wb_clk_i (.I(clknet_3_2__leaf_wb_clk_i),
    .Z(clknet_leaf_16_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_17_wb_clk_i (.I(clknet_3_3__leaf_wb_clk_i),
    .Z(clknet_leaf_17_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_18_wb_clk_i (.I(clknet_3_3__leaf_wb_clk_i),
    .Z(clknet_leaf_18_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_19_wb_clk_i (.I(clknet_opt_2_0_wb_clk_i),
    .Z(clknet_leaf_19_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_20_wb_clk_i (.I(clknet_3_3__leaf_wb_clk_i),
    .Z(clknet_leaf_20_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_21_wb_clk_i (.I(clknet_3_3__leaf_wb_clk_i),
    .Z(clknet_leaf_21_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_22_wb_clk_i (.I(clknet_opt_3_0_wb_clk_i),
    .Z(clknet_leaf_22_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_23_wb_clk_i (.I(clknet_opt_4_0_wb_clk_i),
    .Z(clknet_leaf_23_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_24_wb_clk_i (.I(clknet_3_6__leaf_wb_clk_i),
    .Z(clknet_leaf_24_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_25_wb_clk_i (.I(clknet_3_6__leaf_wb_clk_i),
    .Z(clknet_leaf_25_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_27_wb_clk_i (.I(clknet_3_6__leaf_wb_clk_i),
    .Z(clknet_leaf_27_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_29_wb_clk_i (.I(clknet_3_6__leaf_wb_clk_i),
    .Z(clknet_leaf_29_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_30_wb_clk_i (.I(clknet_3_7__leaf_wb_clk_i),
    .Z(clknet_leaf_30_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_31_wb_clk_i (.I(clknet_3_7__leaf_wb_clk_i),
    .Z(clknet_leaf_31_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_32_wb_clk_i (.I(clknet_3_7__leaf_wb_clk_i),
    .Z(clknet_leaf_32_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_33_wb_clk_i (.I(clknet_3_7__leaf_wb_clk_i),
    .Z(clknet_leaf_33_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_34_wb_clk_i (.I(clknet_3_7__leaf_wb_clk_i),
    .Z(clknet_leaf_34_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_35_wb_clk_i (.I(clknet_3_7__leaf_wb_clk_i),
    .Z(clknet_leaf_35_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_36_wb_clk_i (.I(clknet_3_7__leaf_wb_clk_i),
    .Z(clknet_leaf_36_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_37_wb_clk_i (.I(clknet_3_6__leaf_wb_clk_i),
    .Z(clknet_leaf_37_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_38_wb_clk_i (.I(clknet_3_6__leaf_wb_clk_i),
    .Z(clknet_leaf_38_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_40_wb_clk_i (.I(clknet_3_6__leaf_wb_clk_i),
    .Z(clknet_leaf_40_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_41_wb_clk_i (.I(clknet_3_7__leaf_wb_clk_i),
    .Z(clknet_leaf_41_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_43_wb_clk_i (.I(clknet_3_4__leaf_wb_clk_i),
    .Z(clknet_leaf_43_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_44_wb_clk_i (.I(clknet_3_4__leaf_wb_clk_i),
    .Z(clknet_leaf_44_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_45_wb_clk_i (.I(clknet_3_4__leaf_wb_clk_i),
    .Z(clknet_leaf_45_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_46_wb_clk_i (.I(clknet_3_4__leaf_wb_clk_i),
    .Z(clknet_leaf_46_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_47_wb_clk_i (.I(clknet_3_4__leaf_wb_clk_i),
    .Z(clknet_leaf_47_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_48_wb_clk_i (.I(clknet_3_4__leaf_wb_clk_i),
    .Z(clknet_leaf_48_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_49_wb_clk_i (.I(clknet_3_4__leaf_wb_clk_i),
    .Z(clknet_leaf_49_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_50_wb_clk_i (.I(clknet_3_4__leaf_wb_clk_i),
    .Z(clknet_leaf_50_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_51_wb_clk_i (.I(clknet_3_4__leaf_wb_clk_i),
    .Z(clknet_leaf_51_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_52_wb_clk_i (.I(clknet_3_7__leaf_wb_clk_i),
    .Z(clknet_leaf_52_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_53_wb_clk_i (.I(clknet_3_7__leaf_wb_clk_i),
    .Z(clknet_leaf_53_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_54_wb_clk_i (.I(clknet_3_7__leaf_wb_clk_i),
    .Z(clknet_leaf_54_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_55_wb_clk_i (.I(clknet_3_7__leaf_wb_clk_i),
    .Z(clknet_leaf_55_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_56_wb_clk_i (.I(clknet_3_7__leaf_wb_clk_i),
    .Z(clknet_leaf_56_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_57_wb_clk_i (.I(clknet_3_7__leaf_wb_clk_i),
    .Z(clknet_leaf_57_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_58_wb_clk_i (.I(clknet_3_7__leaf_wb_clk_i),
    .Z(clknet_leaf_58_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_59_wb_clk_i (.I(clknet_3_4__leaf_wb_clk_i),
    .Z(clknet_leaf_59_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_60_wb_clk_i (.I(clknet_3_5__leaf_wb_clk_i),
    .Z(clknet_leaf_60_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_61_wb_clk_i (.I(clknet_3_5__leaf_wb_clk_i),
    .Z(clknet_leaf_61_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_63_wb_clk_i (.I(clknet_3_5__leaf_wb_clk_i),
    .Z(clknet_leaf_63_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_66_wb_clk_i (.I(clknet_3_5__leaf_wb_clk_i),
    .Z(clknet_leaf_66_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_67_wb_clk_i (.I(clknet_3_4__leaf_wb_clk_i),
    .Z(clknet_leaf_67_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_68_wb_clk_i (.I(clknet_3_4__leaf_wb_clk_i),
    .Z(clknet_leaf_68_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_69_wb_clk_i (.I(clknet_3_1__leaf_wb_clk_i),
    .Z(clknet_leaf_69_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_70_wb_clk_i (.I(clknet_3_1__leaf_wb_clk_i),
    .Z(clknet_leaf_70_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_71_wb_clk_i (.I(clknet_3_1__leaf_wb_clk_i),
    .Z(clknet_leaf_71_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_73_wb_clk_i (.I(clknet_3_1__leaf_wb_clk_i),
    .Z(clknet_leaf_73_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_74_wb_clk_i (.I(clknet_3_1__leaf_wb_clk_i),
    .Z(clknet_leaf_74_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_75_wb_clk_i (.I(clknet_3_1__leaf_wb_clk_i),
    .Z(clknet_leaf_75_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_76_wb_clk_i (.I(clknet_3_0__leaf_wb_clk_i),
    .Z(clknet_leaf_76_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_77_wb_clk_i (.I(clknet_3_0__leaf_wb_clk_i),
    .Z(clknet_leaf_77_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_78_wb_clk_i (.I(clknet_3_0__leaf_wb_clk_i),
    .Z(clknet_leaf_78_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_79_wb_clk_i (.I(clknet_3_0__leaf_wb_clk_i),
    .Z(clknet_leaf_79_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_80_wb_clk_i (.I(clknet_3_0__leaf_wb_clk_i),
    .Z(clknet_leaf_80_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_81_wb_clk_i (.I(clknet_3_0__leaf_wb_clk_i),
    .Z(clknet_leaf_81_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_82_wb_clk_i (.I(clknet_3_0__leaf_wb_clk_i),
    .Z(clknet_leaf_82_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_0_wb_clk_i (.I(wb_clk_i),
    .Z(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_0__f_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_1__f_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_2__f_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_3__f_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_4__f_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_5__f_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_6__f_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_7__f_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_opt_1_0_wb_clk_i (.I(clknet_3_3__leaf_wb_clk_i),
    .Z(clknet_opt_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_opt_2_0_wb_clk_i (.I(clknet_3_3__leaf_wb_clk_i),
    .Z(clknet_opt_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_opt_3_0_wb_clk_i (.I(clknet_3_6__leaf_wb_clk_i),
    .Z(clknet_opt_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_opt_4_0_wb_clk_i (.I(clknet_3_6__leaf_wb_clk_i),
    .Z(clknet_opt_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9036__D (.I(_0000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9049__D (.I(_0004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9041__D (.I(_0009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9042__D (.I(_0010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9044__D (.I(_0012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8985__D (.I(_0096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8987__D (.I(_0098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8988__D (.I(_0099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9033__D (.I(_0144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9034__D (.I(_0145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9035__D (.I(_0146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9090__D (.I(_0187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9091__D (.I(_0188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9100__D (.I(_0197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9101__D (.I(_0198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9102__D (.I(_0199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9105__D (.I(_0202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9106__D (.I(_0203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9107__D (.I(_0204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9117__D (.I(_0214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9118__D (.I(_0215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9119__D (.I(_0216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9120__D (.I(_0217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9121__D (.I(_0218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9122__D (.I(_0219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9123__D (.I(_0220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9124__D (.I(_0221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9179__D (.I(_0276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9180__D (.I(_0277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9187__D (.I(_0284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6299__A3 (.I(_0290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4956__I (.I(_0290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4859__A2 (.I(_0290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7228__A3 (.I(_0291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7211__A3 (.I(_0291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4861__A2 (.I(_0291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4960__A2 (.I(_0293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4931__A2 (.I(_0293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4890__A2 (.I(_0293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4862__A2 (.I(_0293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5006__A2 (.I(_0294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4920__B1 (.I(_0294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4863__I (.I(_0294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4881__A2 (.I(_0295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4864__I (.I(_0295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5010__A2 (.I(_0296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4999__A2 (.I(_0296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4886__A2 (.I(_0296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4865__A2 (.I(_0296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5005__A3 (.I(_0298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4957__A2 (.I(_0298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4937__A1 (.I(_0298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4877__A1 (.I(_0298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7907__A1 (.I(_0299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7899__A2 (.I(_0299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5035__A1 (.I(_0299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4869__I (.I(_0299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7975__A1 (.I(_0300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5039__A2 (.I(_0300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5019__A4 (.I(_0300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4877__A2 (.I(_0300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6307__B2 (.I(_0302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5278__A2 (.I(_0302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5135__A2 (.I(_0302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4872__I (.I(_0302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7870__C1 (.I(_0303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5031__A3 (.I(_0303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4985__A2 (.I(_0303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4873__A2 (.I(_0303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7784__C (.I(_0305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7407__A2 (.I(_0305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5078__A1 (.I(_0305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4875__I (.I(_0305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8862__A1 (.I(_0306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7849__B2 (.I(_0306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7664__B2 (.I(_0306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4876__A2 (.I(_0306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4882__A1 (.I(_0308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7902__A1 (.I(_0309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4918__A1 (.I(_0309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4915__A2 (.I(_0309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4880__A1 (.I(_0309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7879__A1 (.I(_0311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4881__B1 (.I(_0311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7594__B (.I(_0314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7540__I (.I(_0314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5232__A1 (.I(_0314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4885__A2 (.I(_0314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7909__A1 (.I(_0315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7863__A2 (.I(_0315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6168__A2 (.I(_0315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4887__A2 (.I(_0315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7236__A1 (.I(_0317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6174__A1 (.I(_0317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5134__A1 (.I(_0317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4889__I (.I(_0317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5490__A1 (.I(_0318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5233__A1 (.I(_0318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4983__A1 (.I(_0318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4890__A1 (.I(_0318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7619__B (.I(_0320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6275__I (.I(_0320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5032__B (.I(_0320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4892__I (.I(_0320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8784__A1 (.I(_0321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7900__A2 (.I(_0321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7275__A2 (.I(_0321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4903__A1 (.I(_0321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7002__C (.I(_0322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6538__C (.I(_0322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4905__I (.I(_0322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4899__A1 (.I(_0322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7053__B (.I(_0323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5128__A2 (.I(_0323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4996__A1 (.I(_0323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4895__I (.I(_0323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7421__I (.I(_0324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7362__A1 (.I(_0324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5490__A3 (.I(_0324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4898__A1 (.I(_0324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7546__B (.I(_0326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7506__I (.I(_0326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7306__I (.I(_0326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4898__A2 (.I(_0326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7906__A2 (.I(_0327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4899__A2 (.I(_0327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7857__A2 (.I(_0330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5229__A1 (.I(_0330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4983__A3 (.I(_0330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4902__A2 (.I(_0330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8428__I (.I(_0333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4984__A1 (.I(_0333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4923__I (.I(_0333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4906__I (.I(_0333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8379__C (.I(_0334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8304__C (.I(_0334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7977__C (.I(_0334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4907__I (.I(_0334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8272__A1 (.I(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7625__A1 (.I(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7478__A1 (.I(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4917__A1 (.I(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7968__A1 (.I(_0336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4927__B2 (.I(_0336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4916__A1 (.I(_0336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4915__A1 (.I(_0336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6485__A1 (.I(_0337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6412__A1 (.I(_0337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5858__A1 (.I(_0337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4910__I (.I(_0337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8030__A2 (.I(_0338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7450__A1 (.I(_0338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7415__I (.I(_0338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4911__I (.I(_0338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7224__B (.I(_0339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6420__A1 (.I(_0339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5038__I (.I(_0339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4912__I (.I(_0339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7711__B2 (.I(_0340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7665__B2 (.I(_0340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7230__A2 (.I(_0340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4916__A2 (.I(_0340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7217__A1 (.I(_0341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5859__A2 (.I(_0341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5851__A1 (.I(_0341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4914__I (.I(_0341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7877__A1 (.I(_0342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6424__A1 (.I(_0342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6416__A1 (.I(_0342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4916__B1 (.I(_0342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4927__A3 (.I(_0343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4916__B2 (.I(_0343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4917__A2 (.I(_0344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7878__A2 (.I(_0345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4920__A3 (.I(_0345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6432__A1 (.I(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6431__A1 (.I(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6412__A2 (.I(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4927__A1 (.I(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8865__C (.I(_0349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8835__C (.I(_0349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8356__C (.I(_0349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4927__A2 (.I(_0349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7788__I (.I(_0350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7575__I (.I(_0350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6347__I (.I(_0350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4925__I (.I(_0350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8813__B (.I(_0351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8621__B (.I(_0351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8610__B (.I(_0351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4926__A2 (.I(_0351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7244__A1 (.I(_0353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7050__A1 (.I(_0353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5032__A1 (.I(_0353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4929__I (.I(_0353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8585__A1 (.I(_0355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8537__A1 (.I(_0355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8519__A1 (.I(_0355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4931__A1 (.I(_0355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8344__B (.I(_0357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7456__A2 (.I(_0357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5020__A1 (.I(_0357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4933__I (.I(_0357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8322__B2 (.I(_0358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7289__A2 (.I(_0358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4992__A3 (.I(_0358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4937__A2 (.I(_0358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7059__I (.I(_0359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5853__A2 (.I(_0359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4964__I (.I(_0359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4935__I (.I(_0359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8787__B1 (.I(_0360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8064__A1 (.I(_0360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7886__I (.I(_0360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4936__A2 (.I(_0360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7870__B1 (.I(_0361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7064__A2 (.I(_0361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4937__A3 (.I(_0361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4958__A2 (.I(_0362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6303__A2 (.I(_0363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4941__A2 (.I(_0363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8838__A2 (.I(_0364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6303__A3 (.I(_0364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6162__A2 (.I(_0364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4940__I (.I(_0364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8593__B1 (.I(_0365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8546__C1 (.I(_0365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5004__I (.I(_0365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4941__A3 (.I(_0365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5011__A1 (.I(_0366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4953__A2 (.I(_0366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6503__A1 (.I(_0367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5863__A2 (.I(_0367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5278__A1 (.I(_0367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4943__I (.I(_0367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8798__A2 (.I(_0368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8479__A2 (.I(_0368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5135__A1 (.I(_0368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4944__I (.I(_0368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7920__B (.I(_0369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6303__A1 (.I(_0369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6109__A2 (.I(_0369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4949__A1 (.I(_0369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5267__A1 (.I(_0370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5220__I (.I(_0370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5110__A1 (.I(_0370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4946__A3 (.I(_0370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6405__A2 (.I(_0371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5058__A2 (.I(_0371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4947__A2 (.I(_0371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6407__A2 (.I(_0373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6282__A1 (.I(_0373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6281__A2 (.I(_0373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4949__A2 (.I(_0373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4953__A3 (.I(_0374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8062__A1 (.I(_0375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4951__I (.I(_0375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7813__A2 (.I(_0377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7740__A2 (.I(_0377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7642__A2 (.I(_0377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4953__B1 (.I(_0377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8579__C (.I(_0380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7899__A3 (.I(_0380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7367__A2 (.I(_0380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4957__A3 (.I(_0380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7901__A1 (.I(_0381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6171__A3 (.I(_0381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5030__A2 (.I(_0381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4957__A4 (.I(_0381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8789__A1 (.I(_0383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6164__A1 (.I(_0383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5031__A1 (.I(_0383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4960__A1 (.I(_0383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7888__A1 (.I(_0385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6178__A1 (.I(_0385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6169__A1 (.I(_0385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4962__I (.I(_0385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7870__A1 (.I(_0386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7709__I (.I(_0386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6344__C (.I(_0386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4963__I (.I(_0386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8872__A1 (.I(_0387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8863__A1 (.I(_0387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7213__A2 (.I(_0387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4978__A1 (.I(_0387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8790__A2 (.I(_0388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8789__C (.I(_0388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8049__B1 (.I(_0388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4965__A1 (.I(_0388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8787__A3 (.I(_0389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7044__A4 (.I(_0389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4977__A2 (.I(_0389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8314__A1 (.I(_0390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7672__A1 (.I(_0390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5848__A2 (.I(_0390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4967__I (.I(_0390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8341__A2 (.I(_0391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8176__A1 (.I(_0391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7655__A1 (.I(_0391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4968__I (.I(_0391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8434__A2 (.I(_0392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8297__A1 (.I(_0392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7995__A2 (.I(_0392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4969__I (.I(_0392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7775__A2 (.I(_0393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7705__A2 (.I(_0393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7522__A2 (.I(_0393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4970__I (.I(_0393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7971__A2 (.I(_0394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7635__A1 (.I(_0394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5019__A2 (.I(_0394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4976__A1 (.I(_0394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8461__A1 (.I(_0395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8395__A1 (.I(_0395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8325__A1 (.I(_0395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4976__A3 (.I(_0395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8248__I (.I(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7284__A2 (.I(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6419__A1 (.I(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4974__I (.I(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8177__C2 (.I(_0398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8143__C2 (.I(_0398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8059__A1 (.I(_0398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4975__I (.I(_0398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8435__B2 (.I(_0399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8365__A1 (.I(_0399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7996__C (.I(_0399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4976__A4 (.I(_0399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4977__B (.I(_0400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4978__A2 (.I(_0401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4993__A2 (.I(_0402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7978__A1 (.I(_0403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4996__A2 (.I(_0403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4980__I (.I(_0403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7662__A1 (.I(_0405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7598__A1 (.I(_0405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7365__B (.I(_0405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4982__I (.I(_0405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7560__A1 (.I(_0406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7509__A1 (.I(_0406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7487__A1 (.I(_0406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4983__A2 (.I(_0406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8342__A1 (.I(_0410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8249__A2 (.I(_0410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6395__A2 (.I(_0410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4987__I (.I(_0410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8361__A2 (.I(_0411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8321__A1 (.I(_0411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7865__A1 (.I(_0411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4988__I (.I(_0411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7634__A2 (.I(_0412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7403__A2 (.I(_0412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6343__B (.I(_0412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4989__I (.I(_0412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6436__A1 (.I(_0413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5039__A1 (.I(_0413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4998__A1 (.I(_0413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4992__A1 (.I(_0413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8068__B (.I(_0414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8029__A1 (.I(_0414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7897__B (.I(_0414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4991__I (.I(_0414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8110__C (.I(_0415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7898__A2 (.I(_0415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5039__B (.I(_0415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4992__A4 (.I(_0415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4993__A4 (.I(_0416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7804__C (.I(_0417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7730__C (.I(_0417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7380__A1 (.I(_0417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4995__I (.I(_0417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7805__A1 (.I(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7771__A1 (.I(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7731__A1 (.I(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4998__A2 (.I(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8494__A1 (.I(_0420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7858__A2 (.I(_0420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4998__B1 (.I(_0420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5000__A2 (.I(_0421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8803__A1 (.I(_0423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7860__A1 (.I(_0423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7775__C (.I(_0423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5002__I (.I(_0423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8822__A1 (.I(_0424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8811__B2 (.I(_0424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8111__C (.I(_0424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5005__A1 (.I(_0424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8417__A1 (.I(_0425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8416__A1 (.I(_0425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7456__A1 (.I(_0425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5005__A2 (.I(_0425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8608__C1 (.I(_0426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8581__A2 (.I(_0426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8565__B1 (.I(_0426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5005__A4 (.I(_0426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5006__B (.I(_0427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8791__B (.I(_0428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5385__A1 (.I(_0428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5051__A1 (.I(_0428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5009__A1 (.I(_0428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8793__C (.I(_0429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7990__A2 (.I(_0429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5017__I (.I(_0429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5009__A2 (.I(_0429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7887__A2 (.I(_0430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5011__A2 (.I(_0430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8877__A1 (.I(_0432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7885__A1 (.I(_0432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5045__I (.I(_0432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5013__I (.I(_0432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7977__A2 (.I(_0433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5086__A1 (.I(_0433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5080__B (.I(_0433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5050__A1 (.I(_0433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7874__A1 (.I(_0434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7455__I (.I(_0434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7048__B (.I(_0434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5015__I (.I(_0434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8445__C (.I(_0435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8285__C (.I(_0435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8158__C (.I(_0435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5016__I (.I(_0435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8396__B (.I(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8103__A1 (.I(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5047__A1 (.I(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5037__A1 (.I(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8212__A1 (.I(_0437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6427__B2 (.I(_0437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6129__A1 (.I(_0437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5019__A1 (.I(_0437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8580__A2 (.I(_0438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7898__C (.I(_0438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5024__A1 (.I(_0438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5019__A3 (.I(_0438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7569__C (.I(_0440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7469__C (.I(_0440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5021__I (.I(_0440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7696__A1 (.I(_0441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7618__A1 (.I(_0441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7516__C (.I(_0441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5037__B1 (.I(_0441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8789__A2 (.I(_0442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7870__A2 (.I(_0442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5859__A3 (.I(_0442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5024__A2 (.I(_0442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5037__B2 (.I(_0444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6302__A1 (.I(_0446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6116__A1 (.I(_0446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5035__B1 (.I(_0446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5030__B1 (.I(_0446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5383__A2 (.I(_0447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5136__A2 (.I(_0447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5028__I (.I(_0447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8606__B (.I(_0448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6310__A2 (.I(_0448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6299__A2 (.I(_0448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5029__A1 (.I(_0448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8791__A1 (.I(_0449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6128__A3 (.I(_0449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5030__B2 (.I(_0449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8838__A1 (.I(_0454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8538__I (.I(_0454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7870__B2 (.I(_0454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5035__B2 (.I(_0454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7573__B2 (.I(_0458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7368__B2 (.I(_0458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7319__B2 (.I(_0458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5050__A2 (.I(_0458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8787__A1 (.I(_0460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7512__I (.I(_0460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5852__A1 (.I(_0460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5041__I (.I(_0460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7693__A2 (.I(_0461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7608__A2 (.I(_0461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7410__A2 (.I(_0461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5044__A1 (.I(_0461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8060__I (.I(_0462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5854__A2 (.I(_0462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5043__I (.I(_0462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8435__A2 (.I(_0463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8252__A2 (.I(_0463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7997__B1 (.I(_0463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5044__A2 (.I(_0463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7976__C (.I(_0465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7229__A1 (.I(_0465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7219__A1 (.I(_0465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5047__B (.I(_0465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8609__A2 (.I(_0466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8594__A2 (.I(_0466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8547__A2 (.I(_0466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5047__C (.I(_0466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8736__A1 (.I(_0468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8707__A1 (.I(_0468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6152__I (.I(_0468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5049__I (.I(_0468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8426__I (.I(_0469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7967__I (.I(_0469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6197__I (.I(_0469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5050__C (.I(_0469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7240__A1 (.I(_0471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5080__A1 (.I(_0471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7970__A1 (.I(_0472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6111__A2 (.I(_0472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5060__A2 (.I(_0472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5055__A1 (.I(_0472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5154__A2 (.I(_0473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5081__A3 (.I(_0473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5066__A3 (.I(_0473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5055__A2 (.I(_0473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5862__I (.I(_0474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5321__A2 (.I(_0474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5055__A3 (.I(_0474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7251__B2 (.I(_0475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6314__A1 (.I(_0475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6313__A2 (.I(_0475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5065__A1 (.I(_0475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6426__A1 (.I(_0476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6323__A1 (.I(_0476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6293__A2 (.I(_0476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5057__A2 (.I(_0476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6394__A1 (.I(_0477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5162__A1 (.I(_0477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5161__A1 (.I(_0477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5059__A1 (.I(_0477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8482__A3 (.I(_0478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5068__A2 (.I(_0478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5059__A3 (.I(_0478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8843__A2 (.I(_0479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5993__A2 (.I(_0479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5878__A2 (.I(_0479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5064__A1 (.I(_0479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8878__A1 (.I(_0480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8706__A1 (.I(_0480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8482__A1 (.I(_0480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5063__A1 (.I(_0480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7217__A3 (.I(_0481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6290__A3 (.I(_0481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5071__I (.I(_0481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5063__A2 (.I(_0481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5328__A2 (.I(_0482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5162__A3 (.I(_0482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5063__A3 (.I(_0482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7250__A1 (.I(_0483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6297__A2 (.I(_0483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5064__A2 (.I(_0483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8868__A1 (.I(_0485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6106__A3 (.I(_0485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5079__A1 (.I(_0485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8876__A1 (.I(_0486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7255__B (.I(_0486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5067__A2 (.I(_0486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6285__A1 (.I(_0487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5079__A2 (.I(_0487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5406__I (.I(_0488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5163__A1 (.I(_0488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5069__I (.I(_0488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8866__A1 (.I(_0489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8559__B2 (.I(_0489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8487__A1 (.I(_0489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5079__A3 (.I(_0489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8787__B2 (.I(_0490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7920__A1 (.I(_0490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6307__A1 (.I(_0490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5078__A2 (.I(_0490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8482__A2 (.I(_0491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7255__A2 (.I(_0491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5162__A2 (.I(_0491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5078__A3 (.I(_0491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5153__A2 (.I(_0492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5148__A2 (.I(_0492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5115__A3 (.I(_0492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5073__I (.I(_0492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8496__A2 (.I(_0493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5385__A2 (.I(_0493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5138__A2 (.I(_0493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5077__A1 (.I(_0493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8891__A1 (.I(_0494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6434__B2 (.I(_0494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5847__A1 (.I(_0494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5075__A1 (.I(_0494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6114__A3 (.I(_0495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5214__A2 (.I(_0495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5076__I (.I(_0495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6316__A3 (.I(_0496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5599__A2 (.I(_0496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5172__A2 (.I(_0496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5077__A2 (.I(_0496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7920__A2 (.I(_0497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5078__A4 (.I(_0497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5080__A2 (.I(_0499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7255__C (.I(_0501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6105__A2 (.I(_0501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5082__I (.I(_0501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8799__A2 (.I(_0502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8588__A2 (.I(_0502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8576__A2 (.I(_0502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5083__I (.I(_0502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8617__A2 (.I(_0503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8524__A2 (.I(_0503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6292__A2 (.I(_0503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5084__B2 (.I(_0503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5086__C (.I(_0505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7056__A2 (.I(_0516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6490__A2 (.I(_0516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5107__A2 (.I(_0516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5137__I (.I(_0518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5109__A2 (.I(_0518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5278__A3 (.I(_0519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5257__A3 (.I(_0519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5135__A3 (.I(_0519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5111__A2 (.I(_0519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8589__B1 (.I(_0520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6730__A2 (.I(_0520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6360__I (.I(_0520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5111__A3 (.I(_0520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5620__I (.I(_0521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5548__C (.I(_0521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5275__I (.I(_0521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5112__I (.I(_0521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5728__A1 (.I(_0523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5693__A2 (.I(_0523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5381__C (.I(_0523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5160__A1 (.I(_0523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6495__A1 (.I(_0524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6486__A1 (.I(_0524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5145__I (.I(_0524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5115__A1 (.I(_0524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5128__A3 (.I(_0525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5116__I (.I(_0525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5490__A4 (.I(_0526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5371__A2 (.I(_0526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5233__A2 (.I(_0526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5127__A2 (.I(_0526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5857__I (.I(_0527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5118__A3 (.I(_0527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5490__A2 (.I(_0529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5128__A1 (.I(_0529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5121__A1 (.I(_0529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7922__A3 (.I(_0530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5133__A3 (.I(_0530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5121__A2 (.I(_0530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7095__I (.I(_0532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5246__I (.I(_0532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5244__A1 (.I(_0532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5124__A1 (.I(_0532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8209__A1 (.I(_0533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7092__I (.I(_0533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5247__A2 (.I(_0533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5124__A2 (.I(_0533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6177__I (.I(_0534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5125__A2 (.I(_0534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6488__A3 (.I(_0536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5371__A3 (.I(_0536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5127__A3 (.I(_0536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5251__I (.I(_0537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5242__I (.I(_0537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5160__A2 (.I(_0537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5345__A2 (.I(_0539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5180__A2 (.I(_0539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5177__I (.I(_0539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5130__I (.I(_0539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7428__I (.I(_0542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7355__I (.I(_0542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5153__A3 (.I(_0542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5133__A2 (.I(_0542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5399__I (.I(_0544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5282__I (.I(_0544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5160__A3 (.I(_0544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5370__I (.I(_0545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5254__I (.I(_0545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5159__A1 (.I(_0545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5385__A3 (.I(_0547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5324__A2 (.I(_0547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5165__A1 (.I(_0547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5138__A4 (.I(_0547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5623__B (.I(_0548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5374__I (.I(_0548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5159__A2 (.I(_0548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6511__A1 (.I(_0549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6376__A1 (.I(_0549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5997__A1 (.I(_0549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5141__A1 (.I(_0549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7233__A1 (.I(_0550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6126__I (.I(_0550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5146__I (.I(_0550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5141__A3 (.I(_0550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8751__A1 (.I(_0551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5331__A1 (.I(_0551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5144__A1 (.I(_0551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7864__A2 (.I(_0552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7049__A3 (.I(_0552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6283__I (.I(_0552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5143__A3 (.I(_0552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8501__B (.I(_0553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6496__A1 (.I(_0553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5144__A2 (.I(_0553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5548__A2 (.I(_0554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5547__A2 (.I(_0554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5159__A3 (.I(_0554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8881__B (.I(_0555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8573__A1 (.I(_0555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6004__A1 (.I(_0555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5158__A1 (.I(_0555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7253__A3 (.I(_0556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7244__B (.I(_0556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5864__A2 (.I(_0556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5149__A2 (.I(_0556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8351__B2 (.I(_0557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7853__A3 (.I(_0557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5149__A3 (.I(_0557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6511__A2 (.I(_0559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5158__A2 (.I(_0559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5993__A3 (.I(_0560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5407__A3 (.I(_0560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5271__A1 (.I(_0560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5157__A1 (.I(_0560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7233__A2 (.I(_0561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5152__I (.I(_0561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7050__A3 (.I(_0562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7037__I (.I(_0562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6104__I (.I(_0562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5155__A2 (.I(_0562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5155__A3 (.I(_0563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6288__A3 (.I(_0564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5155__A4 (.I(_0564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6743__A1 (.I(_0565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5156__I (.I(_0565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8503__A1 (.I(_0566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6502__A1 (.I(_0566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5157__A2 (.I(_0566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5506__I (.I(_0567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5284__I (.I(_0567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5170__I (.I(_0567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5158__B (.I(_0567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5159__A4 (.I(_0568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5728__A4 (.I(_0569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5160__A4 (.I(_0569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8735__A2 (.I(_0570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8706__A2 (.I(_0570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5161__A2 (.I(_0570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5574__A1 (.I(_0571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5426__A1 (.I(_0571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5169__I (.I(_0571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5166__A2 (.I(_0571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8542__A2 (.I(_0572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8491__A4 (.I(_0572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6117__I (.I(_0572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5163__A2 (.I(_0572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8841__B (.I(_0574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8523__B (.I(_0574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8484__B (.I(_0574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5165__A2 (.I(_0574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5574__C (.I(_0576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5426__C (.I(_0576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5335__I (.I(_0576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5167__I (.I(_0576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5666__C (.I(_0582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5531__C (.I(_0582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5226__I (.I(_0582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5173__I (.I(_0582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5773__B2 (.I(_0583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5673__A1 (.I(_0583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5366__B2 (.I(_0583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5228__A1 (.I(_0583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7931__A1 (.I(_0584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5196__A1 (.I(_0584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5183__A1 (.I(_0584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5176__I0 (.I(_0584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6610__A2 (.I(_0589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6562__A1 (.I(_0589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5191__I (.I(_0589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5180__A1 (.I(_0589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5451__A2 (.I(_0592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5219__A1 (.I(_0592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5217__A2 (.I(_0592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5184__A2 (.I(_0592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5657__A2 (.I(_0595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5513__C (.I(_0595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5508__A2 (.I(_0595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5196__A2 (.I(_0595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7916__A1 (.I(_0596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5238__A1 (.I(_0596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5235__I (.I(_0596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5188__A1 (.I(_0596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7913__A1 (.I(_0597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5483__A2 (.I(_0597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5236__A2 (.I(_0597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5188__A2 (.I(_0597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5342__A3 (.I(_0598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5189__I (.I(_0598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6609__A1 (.I(_0601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6607__A1 (.I(_0601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5252__I (.I(_0601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5193__A1 (.I(_0601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5227__A2 (.I(_0605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5219__B (.I(_0605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5217__A1 (.I(_0605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5196__C (.I(_0605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6258__A1 (.I(_0606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5452__A1 (.I(_0606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5197__A2 (.I(_0606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6373__C1 (.I(_0609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5809__I (.I(_0609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5263__A1 (.I(_0609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5201__A1 (.I(_0609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8856__A1 (.I(_0610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8484__A1 (.I(_0610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6373__B2 (.I(_0610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5201__A2 (.I(_0610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5357__A2 (.I(_0611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5202__I (.I(_0611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5810__B (.I(_0612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5263__B (.I(_0612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5207__A2 (.I(_0612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5203__A2 (.I(_0612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5853__A1 (.I(_0614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5210__A1 (.I(_0614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5205__I (.I(_0614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6433__A1 (.I(_0615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6251__A1 (.I(_0615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5599__A1 (.I(_0615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5206__A1 (.I(_0615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5794__B (.I(_0616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5598__I (.I(_0616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5529__A1 (.I(_0616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5207__B (.I(_0616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5452__A2 (.I(_0619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5350__A2 (.I(_0619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5213__A2 (.I(_0619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5212__A2 (.I(_0619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6366__A2 (.I(_0620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5523__I (.I(_0620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5211__I (.I(_0620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6390__A2 (.I(_0621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5455__B (.I(_0621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5352__B (.I(_0621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5212__B (.I(_0621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5449__A1 (.I(_0624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5215__I (.I(_0624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5802__A1 (.I(_0625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5770__A1 (.I(_0625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5600__A1 (.I(_0625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5216__I (.I(_0625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5666__A1 (.I(_0626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5531__A1 (.I(_0626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5224__A1 (.I(_0626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5803__A1 (.I(_0628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5450__B2 (.I(_0628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5361__I (.I(_0628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5224__B2 (.I(_0628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6500__A1 (.I(_0630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5847__A2 (.I(_0630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5256__I (.I(_0630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5221__A2 (.I(_0630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6139__A4 (.I(_0631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5448__A2 (.I(_0631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5364__C (.I(_0631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5222__A2 (.I(_0631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5666__B2 (.I(_0632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5531__B2 (.I(_0632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5450__A1 (.I(_0632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5223__A2 (.I(_0632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5602__A1 (.I(_0636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5431__A1 (.I(_0636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5365__C (.I(_0636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5227__A1 (.I(_0636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8474__A2 (.I(_0638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6534__I0 (.I(_0638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6254__A1 (.I(_0638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5286__A2 (.I(_0638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7488__I (.I(_0639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5232__A2 (.I(_0639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7669__B (.I(_0640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5786__A2 (.I(_0640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5785__A2 (.I(_0640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5231__I (.I(_0640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8504__A2 (.I(_0641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7387__B (.I(_0641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7308__I (.I(_0641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5232__A3 (.I(_0641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5751__A1 (.I(_0643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5234__I (.I(_0643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5748__A1 (.I(_0648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5540__A2 (.I(_0648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5396__B (.I(_0648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5239__A2 (.I(_0648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7309__A2 (.I(_0650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5241__I (.I(_0650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8471__A2 (.I(_0651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7312__A2 (.I(_0651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6532__A1 (.I(_0651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5285__A2 (.I(_0651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5464__A1 (.I(_0654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5391__A2 (.I(_0654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5245__I (.I(_0654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8457__A1 (.I(_0656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5247__A1 (.I(_0656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5464__A2 (.I(_0657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5463__I (.I(_0657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5248__A2 (.I(_0657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7351__A2 (.I(_0659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7350__A2 (.I(_0659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6531__A1 (.I(_0659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5250__I (.I(_0659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8472__A2 (.I(_0660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7305__A1 (.I(_0660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7303__A2 (.I(_0660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5283__A2 (.I(_0660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6687__A1 (.I(_0662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6529__A1 (.I(_0662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6277__A3 (.I(_0662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5253__I (.I(_0662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7924__A1 (.I(_0663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7134__A1 (.I(_0663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5288__I (.I(_0663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5255__A1 (.I(_0663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5745__A2 (.I(_0664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5624__C (.I(_0664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5387__C (.I(_0664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5255__A2 (.I(_0664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8891__A2 (.I(_0666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6436__B2 (.I(_0666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6310__A1 (.I(_0666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5257__A1 (.I(_0666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5471__I (.I(_0667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5258__I (.I(_0667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5829__A1 (.I(_0671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5821__A1 (.I(_0671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5781__A1 (.I(_0671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5262__I (.I(_0671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6364__A2 (.I(_0672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5824__A1 (.I(_0672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5735__I (.I(_0672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5263__A2 (.I(_0672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6527__A1 (.I(_0673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6312__A2 (.I(_0673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5280__A2 (.I(_0673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6790__A1 (.I(_0674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6526__A1 (.I(_0674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6188__I (.I(_0674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5277__A1 (.I(_0674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7351__A1 (.I(_0675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6370__I (.I(_0675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6365__C2 (.I(_0675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5266__I (.I(_0675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7350__A1 (.I(_0676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6521__A1 (.I(_0676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6337__I (.I(_0676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5276__A1 (.I(_0676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8791__C (.I(_0677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6300__I (.I(_0677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5268__A2 (.I(_0677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8619__A2 (.I(_0678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5270__A2 (.I(_0678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8212__A2 (.I(_0679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7887__A3 (.I(_0679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5270__A3 (.I(_0679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5273__I (.I(_0681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5272__I (.I(_0681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5470__I (.I(_0688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5279__I (.I(_0688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5774__A1 (.I(_0694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5559__C (.I(_0694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5339__I (.I(_0694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5285__C (.I(_0694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8739__A1 (.I(_0696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8710__A1 (.I(_0696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5287__I (.I(_0696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5336__A2 (.I(_0697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8514__A1 (.I(_0698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6183__A1 (.I(_0698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5881__A1 (.I(_0698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5325__I0 (.I(_0698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8010__A1 (.I(_0699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6386__A1 (.I(_0699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6226__A1 (.I(_0699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5290__I (.I(_0699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8481__A1 (.I(_0700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6438__A1 (.I(_0700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5960__I (.I(_0700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5293__A1 (.I(_0700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8523__A1 (.I(_0702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7102__A2 (.I(_0702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5307__A2 (.I(_0702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5293__A2 (.I(_0702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5704__A2 (.I(_0704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5568__A2 (.I(_0704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5419__B1 (.I(_0704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5295__I (.I(_0704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5939__A2 (.I(_0705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5722__A2 (.I(_0705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5720__A2 (.I(_0705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5306__A2 (.I(_0705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6387__A1 (.I(_0708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6226__A2 (.I(_0708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5962__I (.I(_0708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5299__A2 (.I(_0708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5704__B1 (.I(_0710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5634__B1 (.I(_0710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5568__B1 (.I(_0710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5301__I (.I(_0710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6972__A2 (.I(_0711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5722__B1 (.I(_0711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5720__B1 (.I(_0711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5306__B1 (.I(_0711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5568__C2 (.I(_0713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5497__A2 (.I(_0713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5412__I (.I(_0713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5304__I (.I(_0713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8760__A2 (.I(_0715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5567__A2 (.I(_0715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5319__A2 (.I(_0715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5306__C2 (.I(_0715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5638__I (.I(_0717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5413__I (.I(_0717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5308__I (.I(_0717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5706__B1 (.I(_0718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5565__C1 (.I(_0718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5421__B1 (.I(_0718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5309__I (.I(_0718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5869__A2 (.I(_0719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5570__A2 (.I(_0719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5319__B1 (.I(_0719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5314__A2 (.I(_0719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8200__C (.I(_0721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5640__I (.I(_0721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5416__I (.I(_0721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5312__I (.I(_0721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8262__C (.I(_0722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8075__C (.I(_0722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5422__I (.I(_0722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5313__I (.I(_0722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8811__A2 (.I(_0723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8282__B2 (.I(_0723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5320__B2 (.I(_0723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5314__B (.I(_0723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5636__A2 (.I(_0725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5565__A2 (.I(_0725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5495__A2 (.I(_0725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5317__A2 (.I(_0725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5565__B1 (.I(_0726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5495__B1 (.I(_0726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5417__B1 (.I(_0726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5317__B1 (.I(_0726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8327__A2 (.I(_0730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7135__A1 (.I(_0730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5325__I1 (.I(_0730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7257__A1 (.I(_0731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6305__A2 (.I(_0731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6105__A1 (.I(_0731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5322__I (.I(_0731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8816__B (.I(_0732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8588__B2 (.I(_0732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7132__I (.I(_0732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5323__I (.I(_0732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8809__A1 (.I(_0733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8808__C (.I(_0733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8617__B2 (.I(_0733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5324__A1 (.I(_0733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6418__A1 (.I(_0736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6291__A1 (.I(_0736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6115__B (.I(_0736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5327__I (.I(_0736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8208__A1 (.I(_0737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7129__I (.I(_0737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6118__I (.I(_0737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5330__A1 (.I(_0737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6291__A2 (.I(_0738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6106__A2 (.I(_0738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5329__I (.I(_0738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8797__A2 (.I(_0739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7243__A1 (.I(_0739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6120__A1 (.I(_0739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5330__A2 (.I(_0739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8751__A2 (.I(_0740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6899__A1 (.I(_0740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6536__A1 (.I(_0740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5331__A2 (.I(_0740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8725__I (.I(_0741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8704__I (.I(_0741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5332__A2 (.I(_0741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5453__A1 (.I(_0750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5366__B1 (.I(_0750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5348__A1 (.I(_0750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6593__A2 (.I(_0752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6549__B2 (.I(_0752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5367__I (.I(_0752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5344__I (.I(_0752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6739__A1 (.I(_0753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5888__I0 (.I(_0753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5410__A1 (.I(_0753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5345__A1 (.I(_0753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5346__B2 (.I(_0754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5356__A2 (.I(_0755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5347__I (.I(_0755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6272__A2 (.I(_0758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5365__A2 (.I(_0758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5353__A1 (.I(_0758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5352__A1 (.I(_0758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5363__A1 (.I(_0764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5362__A1 (.I(_0764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5356__A1 (.I(_0764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5771__A1 (.I(_0770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5601__A1 (.I(_0770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5521__A1 (.I(_0770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5365__A1 (.I(_0770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8519__A2 (.I(_0775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6744__A1 (.I(_0775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6253__A1 (.I(_0775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5402__A2 (.I(_0775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6750__A1 (.I(_0777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6608__A1 (.I(_0777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6277__A2 (.I(_0777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5369__I (.I(_0777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8817__A1 (.I(_0778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7007__A1 (.I(_0778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6187__I (.I(_0778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5388__A1 (.I(_0778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5696__A2 (.I(_0779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5695__B (.I(_0779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5625__A2 (.I(_0779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5388__A2 (.I(_0779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5610__I (.I(_0780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5556__A1 (.I(_0780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5372__I (.I(_0780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5826__A1 (.I(_0781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5747__A1 (.I(_0781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5746__B (.I(_0781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5388__B (.I(_0781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6737__A1 (.I(_0782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6180__I (.I(_0782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5810__A2 (.I(_0782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5387__A1 (.I(_0782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5695__A2 (.I(_0783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5624__A2 (.I(_0783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5387__A2 (.I(_0783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5386__B (.I(_0783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8052__A1 (.I(_0784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7377__A2 (.I(_0784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6374__I (.I(_0784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5376__I (.I(_0784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7390__A1 (.I(_0786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6734__A1 (.I(_0786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6368__B2 (.I(_0786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5378__I (.I(_0786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8063__A1 (.I(_0787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8055__A1 (.I(_0787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6338__I (.I(_0787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5381__A1 (.I(_0787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5692__A2 (.I(_0788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5621__A2 (.I(_0788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5381__A2 (.I(_0788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5380__A2 (.I(_0788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8563__A1 (.I(_0791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8546__C2 (.I(_0791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6736__A1 (.I(_0791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5386__A1 (.I(_0791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8578__B1 (.I(_0793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6332__A1 (.I(_0793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6326__B (.I(_0793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5385__A4 (.I(_0793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5623__A2 (.I(_0794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5386__A2 (.I(_0794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5535__C (.I(_0798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5397__A2 (.I(_0798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5392__A2 (.I(_0798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5391__A1 (.I(_0798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5732__A1 (.I(_0799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5553__A2 (.I(_0799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5391__B (.I(_0799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8518__A2 (.I(_0802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7390__A2 (.I(_0802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6740__A1 (.I(_0802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5394__A2 (.I(_0802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5608__B2 (.I(_0804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5604__A1 (.I(_0804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5534__I (.I(_0804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5396__A2 (.I(_0804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8516__A2 (.I(_0806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7382__A2 (.I(_0806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7356__A2 (.I(_0806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5398__I (.I(_0806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6742__A1 (.I(_0807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5400__B1 (.I(_0807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5728__A3 (.I(_0808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5631__C (.I(_0808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5559__A1 (.I(_0808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5400__B2 (.I(_0808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8742__A1 (.I(_0811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8715__B2 (.I(_0811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5426__A2 (.I(_0811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8044__B (.I(_0812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7208__I (.I(_0812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6123__I (.I(_0812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5404__I (.I(_0812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8284__C (.I(_0813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7272__A1 (.I(_0813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6316__A1 (.I(_0813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5405__I (.I(_0813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8065__B (.I(_0814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7997__C (.I(_0814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6108__I (.I(_0814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5407__A1 (.I(_0814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8601__A1 (.I(_0815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8544__A1 (.I(_0815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7130__A2 (.I(_0815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5407__A2 (.I(_0815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5411__I (.I(_0816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5408__I (.I(_0816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5706__A2 (.I(_0821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5496__A2 (.I(_0821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5494__A2 (.I(_0821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5414__A2 (.I(_0821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5636__B1 (.I(_0822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5496__B1 (.I(_0822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5494__B1 (.I(_0822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5414__B1 (.I(_0822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5708__A2 (.I(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5642__A2 (.I(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5499__A2 (.I(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5417__A2 (.I(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8155__C (.I(_0825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5708__C (.I(_0825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5495__C (.I(_0825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5417__C (.I(_0825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5708__B1 (.I(_0827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5642__B1 (.I(_0827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5499__B1 (.I(_0827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5421__A2 (.I(_0827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8156__A1 (.I(_0831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5709__A1 (.I(_0831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5643__A1 (.I(_0831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5423__B2 (.I(_0831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8353__A2 (.I(_0832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7147__A1 (.I(_0832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5424__A2 (.I(_0832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5525__A1 (.I(_0838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5431__A2 (.I(_0838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5659__A2 (.I(_0840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5658__A2 (.I(_0840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5439__A2 (.I(_0840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5434__A2 (.I(_0840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5893__I0 (.I(_0845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5502__A1 (.I(_0845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5438__A1 (.I(_0845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5525__A2 (.I(_0847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5441__A2 (.I(_0847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5440__A2 (.I(_0847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6259__A1 (.I(_0848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5519__A3 (.I(_0848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5449__A2 (.I(_0848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5442__A1 (.I(_0848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5596__A1 (.I(_0849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5445__I (.I(_0849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5442__A2 (.I(_0849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6259__A2 (.I(_0853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5529__A2 (.I(_0853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5520__A1 (.I(_0853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5450__A2 (.I(_0853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6125__A2 (.I(_0855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5667__A1 (.I(_0855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5448__A3 (.I(_0855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5802__C (.I(_0856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5600__C (.I(_0856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5507__I (.I(_0856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5449__B (.I(_0856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6796__A1 (.I(_0866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5493__I0 (.I(_0866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5485__A2 (.I(_0870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5466__B1 (.I(_0870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8535__A2 (.I(_0874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7431__A2 (.I(_0874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7392__A2 (.I(_0874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5467__I (.I(_0874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7393__A2 (.I(_0875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6792__A1 (.I(_0875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5482__A2 (.I(_0875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6612__B2 (.I(_0876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6590__A1 (.I(_0876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6277__A1 (.I(_0876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5469__I (.I(_0876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8807__A1 (.I(_0877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6791__A1 (.I(_0877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6193__I (.I(_0877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5481__A1 (.I(_0877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6890__A1 (.I(_0880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6199__I (.I(_0880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5624__A1 (.I(_0880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5478__A1 (.I(_0880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8134__A1 (.I(_0881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7431__A1 (.I(_0881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6378__I (.I(_0881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5474__I (.I(_0881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7392__A1 (.I(_0882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6786__A1 (.I(_0882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6365__A1 (.I(_0882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5475__I (.I(_0882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7385__A1 (.I(_0883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7381__I (.I(_0883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6339__I (.I(_0883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5477__A1 (.I(_0883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5829__B2 (.I(_0892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5679__A3 (.I(_0892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5608__C2 (.I(_0892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5485__A1 (.I(_0892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7424__A2 (.I(_0893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7384__A1 (.I(_0893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5488__A1 (.I(_0893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7424__A3 (.I(_0895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7384__A2 (.I(_0895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5488__A2 (.I(_0895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8536__A2 (.I(_0896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7385__A2 (.I(_0896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6794__A1 (.I(_0896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5492__I1 (.I(_0896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5832__A1 (.I(_0899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5747__C (.I(_0899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5492__S (.I(_0899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8745__A1 (.I(_0901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8718__B2 (.I(_0901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5503__A2 (.I(_0901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8185__C (.I(_0905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8115__C (.I(_0905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5566__I (.I(_0905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5498__I (.I(_0905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8073__C (.I(_0906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8022__B (.I(_0906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5569__A1 (.I(_0906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5499__C (.I(_0906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8376__A2 (.I(_0908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7153__A1 (.I(_0908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5501__A2 (.I(_0908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8855__A2 (.I(_0914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5805__A1 (.I(_0914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5770__C (.I(_0914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5533__A1 (.I(_0914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5533__A2 (.I(_0916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5530__A1 (.I(_0916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5516__A1 (.I(_0916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5515__A1 (.I(_0916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6807__A1 (.I(_0918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6574__A1 (.I(_0918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5542__I (.I(_0918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5512__A1 (.I(_0918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5596__A3 (.I(_0926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5529__A4 (.I(_0926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5520__A2 (.I(_0926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5804__A1 (.I(_0930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5764__B (.I(_0930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5594__B (.I(_0930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5524__I (.I(_0930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8861__A1 (.I(_0931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8854__A1 (.I(_0931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5671__A1 (.I(_0931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5532__A1 (.I(_0931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8850__A2 (.I(_0934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5593__A2 (.I(_0934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5528__A2 (.I(_0934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8553__A2 (.I(_0940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6839__A1 (.I(_0940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6254__A2 (.I(_0940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5560__A2 (.I(_0940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5828__A1 (.I(_0941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5749__B2 (.I(_0941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5680__B2 (.I(_0941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5537__A1 (.I(_0941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5554__B1 (.I(_0943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5537__A2 (.I(_0943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5607__A2 (.I(_0945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5553__A1 (.I(_0945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5540__A1 (.I(_0945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8552__A2 (.I(_0948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6838__A1 (.I(_0948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5559__A2 (.I(_0948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6835__A1 (.I(_0949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6278__A4 (.I(_0949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5562__I (.I(_0949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5551__A1 (.I(_0949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8526__B2 (.I(_0950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6834__A1 (.I(_0950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6194__A1 (.I(_0950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5550__A1 (.I(_0950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6830__I (.I(_0951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5678__A1 (.I(_0951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5627__A1 (.I(_0951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5549__A1 (.I(_0951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8132__A1 (.I(_0952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8131__A1 (.I(_0952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7444__A2 (.I(_0952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5546__I (.I(_0952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7499__A1 (.I(_0953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6831__A1 (.I(_0953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6340__I (.I(_0953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5547__A1 (.I(_0953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5549__B (.I(_0955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7499__A2 (.I(_0961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7498__A2 (.I(_0961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5555__I (.I(_0961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8551__A2 (.I(_0962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7434__A2 (.I(_0962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6837__A1 (.I(_0962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5556__A2 (.I(_0962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8749__A1 (.I(_0967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8721__A1 (.I(_0967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5561__I (.I(_0967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8567__A1 (.I(_0969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7159__B2 (.I(_0969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6201__A1 (.I(_0969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5563__I (.I(_0969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7945__A1 (.I(_0970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5900__I0 (.I(_0970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5564__A1 (.I(_0970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5571__A1 (.I(_0972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8809__A2 (.I(_0973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8023__A1 (.I(_0973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5723__C (.I(_0973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5567__B (.I(_0973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8397__A2 (.I(_0978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7158__A1 (.I(_0978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5572__A2 (.I(_0978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5840__A2 (.I(_0983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5778__A2 (.I(_0983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5714__A2 (.I(_0983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5648__A2 (.I(_0983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6843__A1 (.I(_0988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6647__A1 (.I(_0988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5611__I (.I(_0988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5583__A1 (.I(_0988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6257__A1 (.I(_0995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5669__A1 (.I(_0995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5597__A1 (.I(_0995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5590__I (.I(_0995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5669__A2 (.I(_0999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5595__A2 (.I(_0999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5594__A2 (.I(_0999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8853__C (.I(_1004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5768__A1 (.I(_1004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5672__A1 (.I(_1004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5601__B2 (.I(_1004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5802__B2 (.I(_1005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5770__B2 (.I(_1005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5600__B2 (.I(_1005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8572__A2 (.I(_1009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6886__A1 (.I(_1009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6255__A1 (.I(_1009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5633__A2 (.I(_1009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5628__A2 (.I(_1012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5608__B1 (.I(_1012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7492__A2 (.I(_1014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5609__I (.I(_1014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8571__A2 (.I(_1015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7548__A2 (.I(_1015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6894__A1 (.I(_1015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5632__A2 (.I(_1015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6891__A1 (.I(_1017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6879__A1 (.I(_1017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6278__A3 (.I(_1017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5612__I (.I(_1017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7951__A1 (.I(_1018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5905__I (.I(_1018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5645__A1 (.I(_1018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5625__A1 (.I(_1018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8219__A1 (.I(_1019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8218__A1 (.I(_1019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7492__A1 (.I(_1019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5614__I (.I(_1019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7536__A2 (.I(_1021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6388__A2 (.I(_1021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6376__A2 (.I(_1021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5616__I (.I(_1021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8171__A1 (.I(_1022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6887__A1 (.I(_1022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6364__C2 (.I(_1022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5617__I (.I(_1022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8177__A1 (.I(_1023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7501__A1 (.I(_1023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6333__I (.I(_1023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5621__A1 (.I(_1023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8607__A1 (.I(_1028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8593__B2 (.I(_1028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5744__A1 (.I(_1028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5623__A1 (.I(_1028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5624__B2 (.I(_1029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7543__A2 (.I(_1034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7542__A2 (.I(_1034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5629__I (.I(_1034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8570__A2 (.I(_1035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7501__A2 (.I(_1035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6893__A1 (.I(_1035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5630__A2 (.I(_1035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8750__A1 (.I(_1039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8723__B2 (.I(_1039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5647__A2 (.I(_1039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5723__A2 (.I(_1043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5721__A2 (.I(_1043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5707__A2 (.I(_1043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5639__A2 (.I(_1043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5723__B1 (.I(_1044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5721__B1 (.I(_1044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5707__B1 (.I(_1044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5639__B1 (.I(_1044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8204__B2 (.I(_1046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8183__C (.I(_1046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8118__C (.I(_1046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5641__I (.I(_1046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8278__C (.I(_1047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8266__B2 (.I(_1047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5721__C (.I(_1047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5642__C (.I(_1047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8423__A2 (.I(_1049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7164__A1 (.I(_1049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5644__A2 (.I(_1049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6212__I (.I(_1055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5698__A1 (.I(_1055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5680__A1 (.I(_1055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5654__A1 (.I(_1055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7955__I1 (.I(_1056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5664__A1 (.I(_1056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5659__A1 (.I(_1056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5653__A1 (.I(_1056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5781__A2 (.I(_1057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5780__A2 (.I(_1057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5757__A2 (.I(_1057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5653__A2 (.I(_1057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8585__A2 (.I(_1078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6909__A1 (.I(_1078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6255__A2 (.I(_1078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5703__A2 (.I(_1078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5820__A2 (.I(_1079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5730__A2 (.I(_1079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5676__A1 (.I(_1079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5731__A1 (.I(_1082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5697__A1 (.I(_1082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5679__A1 (.I(_1082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5697__A2 (.I(_1083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5679__A2 (.I(_1083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7589__A2 (.I(_1085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7588__A2 (.I(_1085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5681__I (.I(_1085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8584__A2 (.I(_1086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7550__A2 (.I(_1086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6908__A1 (.I(_1086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5702__A2 (.I(_1086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6905__A1 (.I(_1087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6867__A1 (.I(_1087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6278__A2 (.I(_1087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5683__I (.I(_1087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6137__A1 (.I(_1088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5915__I (.I(_1088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5711__A1 (.I(_1088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5696__A1 (.I(_1088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6957__A1 (.I(_1089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6365__B1 (.I(_1089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5818__A1 (.I(_1089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5685__I (.I(_1089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8608__C2 (.I(_1090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6326__A1 (.I(_1090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6217__A1 (.I(_1090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5693__A1 (.I(_1090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7602__B1 (.I(_1091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7562__A2 (.I(_1091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7535__A2 (.I(_1091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5687__I (.I(_1091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8239__A1 (.I(_1092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8238__A1 (.I(_1092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7589__A1 (.I(_1092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5688__I (.I(_1092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7550__A1 (.I(_1094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6901__A1 (.I(_1094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6364__B2 (.I(_1094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5690__I (.I(_1094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8222__A1 (.I(_1095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6336__A2 (.I(_1095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6135__I (.I(_1095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5692__A1 (.I(_1095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6904__A1 (.I(_1099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6328__A2 (.I(_1099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6207__A1 (.I(_1099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5695__A1 (.I(_1099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7581__A2 (.I(_1103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7580__A2 (.I(_1103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5699__I (.I(_1103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8583__A2 (.I(_1104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7545__A2 (.I(_1104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6900__I (.I(_1104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5700__A2 (.I(_1104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8752__A1 (.I(_1108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8728__A1 (.I(_1108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5713__A2 (.I(_1108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8446__A2 (.I(_1114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7169__A1 (.I(_1114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5710__A2 (.I(_1114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6919__A1 (.I(_1120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6751__A1 (.I(_1120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6278__A1 (.I(_1120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5717__I (.I(_1120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6933__A1 (.I(_1121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5923__I (.I(_1121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5745__A1 (.I(_1121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5718__I (.I(_1121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7960__A1 (.I(_1122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6313__A1 (.I(_1122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5719__A1 (.I(_1122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8462__A2 (.I(_1128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7175__A1 (.I(_1128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5725__A2 (.I(_1128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7125__A1 (.I(_1131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6121__A1 (.I(_1131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5863__A1 (.I(_1131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5729__A1 (.I(_1131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8734__A2 (.I(_1132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8703__A2 (.I(_1132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5729__A2 (.I(_1132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7579__A2 (.I(_1137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5734__I (.I(_1137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8598__A2 (.I(_1138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7653__A2 (.I(_1138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6927__I (.I(_1138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5747__A2 (.I(_1138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8847__A1 (.I(_1139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8619__B2 (.I(_1139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6222__A1 (.I(_1139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5743__A1 (.I(_1139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8252__A1 (.I(_1143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6365__B2 (.I(_1143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6334__I (.I(_1143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5742__A1 (.I(_1143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6928__A1 (.I(_1144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5741__A1 (.I(_1144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7587__A2 (.I(_1153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5750__I (.I(_1153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8599__A2 (.I(_1154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7646__A2 (.I(_1154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6935__A1 (.I(_1154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5751__A2 (.I(_1154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8600__A2 (.I(_1177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6936__I0 (.I(_1177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6255__A3 (.I(_1177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5774__A2 (.I(_1177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8756__A1 (.I(_1179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8731__A1 (.I(_1179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5776__A2 (.I(_1179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5777__C (.I(_1180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6916__A1 (.I(_1186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6851__A1 (.I(_1186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6802__A1 (.I(_1186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5784__I (.I(_1186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6945__A1 (.I(_1187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6944__A1 (.I(_1187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5807__I (.I(_1187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5786__A1 (.I(_1187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8853__A2 (.I(_1196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5795__A2 (.I(_1196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5794__A2 (.I(_1196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8614__A2 (.I(_1209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6962__A1 (.I(_1209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6274__A2 (.I(_1209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5835__A2 (.I(_1209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6958__A1 (.I(_1210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6399__A1 (.I(_1210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6279__B (.I(_1210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5808__I (.I(_1210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7180__A1 (.I(_1211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5935__A1 (.I(_1211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5837__I (.I(_1211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5819__A1 (.I(_1211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8885__B (.I(_1212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8842__A1 (.I(_1212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8558__A1 (.I(_1212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5810__A1 (.I(_1212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6956__A1 (.I(_1213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6361__B2 (.I(_1213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6332__A2 (.I(_1213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5817__A2 (.I(_1213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6953__I (.I(_1214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6387__C2 (.I(_1214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6373__A2 (.I(_1214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5812__I (.I(_1214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7668__A1 (.I(_1215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7276__I (.I(_1215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6418__A2 (.I(_1215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5813__I (.I(_1215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8142__A2 (.I(_1216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7649__A1 (.I(_1216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7098__I (.I(_1216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5816__A1 (.I(_1216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8620__A1 (.I(_1217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7991__A1 (.I(_1217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6955__A1 (.I(_1217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5815__A1 (.I(_1217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6282__B2 (.I(_1225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5823__A2 (.I(_1225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7673__A2 (.I(_1227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7672__A2 (.I(_1227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5825__I (.I(_1227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8612__A2 (.I(_1228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7655__A2 (.I(_1228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6960__A1 (.I(_1228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5826__A2 (.I(_1228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7669__A2 (.I(_1233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7668__A2 (.I(_1233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5831__I (.I(_1233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8613__A2 (.I(_1234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7649__A2 (.I(_1234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6961__A1 (.I(_1234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5832__A2 (.I(_1234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8759__A1 (.I(_1238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8733__A1 (.I(_1238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5836__A2 (.I(_1238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8621__A1 (.I(_1240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7976__A1 (.I(_1240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6223__A1 (.I(_1240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5838__A1 (.I(_1240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5840__B2 (.I(_1242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7045__A3 (.I(_1244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5843__I (.I(_1244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7043__I (.I(_1245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6429__A2 (.I(_1245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5855__A1 (.I(_1245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5853__B1 (.I(_1245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7216__I (.I(_1246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5850__A2 (.I(_1246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5845__A1 (.I(_1246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7855__A2 (.I(_1247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7238__I (.I(_1247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5876__A2 (.I(_1247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5846__A2 (.I(_1247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8799__A3 (.I(_1248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8502__C (.I(_1248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6161__A3 (.I(_1248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5849__A2 (.I(_1248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8794__A2 (.I(_1249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5860__A2 (.I(_1249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5852__A2 (.I(_1249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5849__A3 (.I(_1249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7877__A3 (.I(_1252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7871__B2 (.I(_1252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7269__A1 (.I(_1252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5851__A2 (.I(_1252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7246__A3 (.I(_1253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7227__A2 (.I(_1253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7225__I (.I(_1253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5854__A3 (.I(_1253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5854__A4 (.I(_1255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5855__B (.I(_1256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8794__B2 (.I(_1258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8793__A2 (.I(_1258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7887__A1 (.I(_1258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5861__A2 (.I(_1258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8001__A2 (.I(_1259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7919__I (.I(_1259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7411__C (.I(_1259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5858__A3 (.I(_1259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6508__A2 (.I(_1260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5860__A3 (.I(_1260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5860__A4 (.I(_1261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5866__B (.I(_1263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8798__A3 (.I(_1264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8479__A3 (.I(_1264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6109__A3 (.I(_1264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5863__A3 (.I(_1264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7980__A2 (.I(_1266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7251__A2 (.I(_1266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7240__A2 (.I(_1266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5865__A3 (.I(_1266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6004__A2 (.I(_1267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5908__I (.I(_1267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5871__I (.I(_1267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5866__C (.I(_1267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6458__I (.I(_1268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5989__I (.I(_1268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5867__I (.I(_1268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5912__I (.I(_1271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5904__I (.I(_1271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5883__I (.I(_1271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5870__I (.I(_1271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8126__A3 (.I(_1274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8047__A1 (.I(_1274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7329__A1 (.I(_1274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5873__I (.I(_1274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8086__A2 (.I(_1275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8042__A2 (.I(_1275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7990__A1 (.I(_1275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5874__I (.I(_1275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7995__A1 (.I(_1276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7989__I (.I(_1276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7279__A1 (.I(_1276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5875__I (.I(_1276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8031__A1 (.I(_1277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8007__B2 (.I(_1277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7267__I (.I(_1277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5880__A1 (.I(_1277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7250__A2 (.I(_1278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7249__A2 (.I(_1278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7241__A2 (.I(_1278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5877__I (.I(_1278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7966__A3 (.I(_1279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7256__A1 (.I(_1279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7243__A2 (.I(_1279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5878__A3 (.I(_1279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5997__A2 (.I(_1280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5927__A2 (.I(_1280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5879__I (.I(_1280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6970__I (.I(_1283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5882__I (.I(_1283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6070__A1 (.I(_1284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5971__A1 (.I(_1284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5943__A1 (.I(_1284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5885__A2 (.I(_1284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8104__A1 (.I(_1287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8058__A1 (.I(_1287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8042__A1 (.I(_1287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5887__I (.I(_1287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8084__A1 (.I(_1288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7367__A1 (.I(_1288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7339__B (.I(_1288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5888__I1 (.I(_1288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6072__A1 (.I(_1290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5973__A1 (.I(_1290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5945__A1 (.I(_1290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5891__A2 (.I(_1290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7447__A1 (.I(_1292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7416__A1 (.I(_1292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5893__I1 (.I(_1292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6980__I (.I(_1293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5894__I (.I(_1293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6074__A1 (.I(_1294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5975__A1 (.I(_1294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5947__A1 (.I(_1294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5896__A2 (.I(_1294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8214__A3 (.I(_1296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8195__A2 (.I(_1296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7445__A1 (.I(_1296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5898__I (.I(_1296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8167__A1 (.I(_1297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8164__A1 (.I(_1297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8142__A1 (.I(_1297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5899__I (.I(_1297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8163__A1 (.I(_1298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8127__A1 (.I(_1298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7473__A1 (.I(_1298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5900__I1 (.I(_1298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6983__I (.I(_1299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5901__I (.I(_1299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6076__A1 (.I(_1300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5977__A1 (.I(_1300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5949__A1 (.I(_1300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5903__A2 (.I(_1300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8569__A1 (.I(_1303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7165__B2 (.I(_1303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6208__A1 (.I(_1303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5910__A1 (.I(_1303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8214__A2 (.I(_1304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8195__A1 (.I(_1304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7479__A1 (.I(_1304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5907__I (.I(_1304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8193__A1 (.I(_1305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8168__A1 (.I(_1305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7527__A1 (.I(_1305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5909__A1 (.I(_1305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6986__I (.I(_1308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5911__I (.I(_1308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6080__A1 (.I(_1309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5981__A1 (.I(_1309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5953__A1 (.I(_1309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5914__A2 (.I(_1309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5937__A2 (.I(_1310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5930__A2 (.I(_1310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5921__A2 (.I(_1310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5913__A2 (.I(_1310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8596__A1 (.I(_1312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7170__B2 (.I(_1312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6214__A1 (.I(_1312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5919__A1 (.I(_1312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8214__A1 (.I(_1313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7603__A1 (.I(_1313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7535__A1 (.I(_1313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5917__I (.I(_1313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8232__A1 (.I(_1314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8206__A1 (.I(_1314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7571__A1 (.I(_1314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5918__A1 (.I(_1314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6991__I (.I(_1316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5920__I (.I(_1316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6082__A1 (.I(_1317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5983__A1 (.I(_1317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5955__A1 (.I(_1317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5922__A2 (.I(_1317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8610__A1 (.I(_1319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7176__B2 (.I(_1319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6218__A1 (.I(_1319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5928__A1 (.I(_1319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8249__A1 (.I(_1321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8247__A1 (.I(_1321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8234__A1 (.I(_1321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5926__I (.I(_1321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8271__A1 (.I(_1322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7622__A1 (.I(_1322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7619__A1 (.I(_1322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5927__A1 (.I(_1322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6994__I (.I(_1324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5929__I (.I(_1324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6084__A1 (.I(_1325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5985__A1 (.I(_1325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5957__A1 (.I(_1325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5931__A2 (.I(_1325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8304__A1 (.I(_1328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8288__A1 (.I(_1328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8284__A1 (.I(_1328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5934__A1 (.I(_1328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6997__I (.I(_1330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5936__I (.I(_1330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6086__A1 (.I(_1331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5987__A1 (.I(_1331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5959__A1 (.I(_1331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5938__A2 (.I(_1331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5951__I (.I(_1333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5950__I (.I(_1333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5941__I (.I(_1333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5940__I (.I(_1333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5948__A2 (.I(_1335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5946__A2 (.I(_1335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5944__A2 (.I(_1335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5942__A2 (.I(_1335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8825__I0 (.I(_1349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8663__A2 (.I(_1349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8623__A2 (.I(_1349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5966__A1 (.I(_1349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8806__A1 (.I(_1350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8541__A1 (.I(_1350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5988__I (.I(_1350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5965__I (.I(_1350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5979__I (.I(_1353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5978__I (.I(_1353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5969__I (.I(_1353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5968__I (.I(_1353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6020__I (.I(_1368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5991__I (.I(_1368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6063__A2 (.I(_1369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6055__A2 (.I(_1369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6009__I (.I(_1369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5992__I (.I(_1369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6041__A1 (.I(_1370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6030__A1 (.I(_1370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6022__A1 (.I(_1370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6011__A1 (.I(_1370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6015__I (.I(_1371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5994__I (.I(_1371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6043__A2 (.I(_1375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6025__A2 (.I(_1375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6014__I (.I(_1375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5998__I (.I(_1375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8357__A2 (.I(_1378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7766__A2 (.I(_1378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7716__A1 (.I(_1378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6001__I (.I(_1378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8334__A1 (.I(_1381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7711__A1 (.I(_1381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7708__A1 (.I(_1381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6005__A1 (.I(_1381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6006__A3 (.I(_1383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6457__I (.I(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6008__I (.I(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6064__A1 (.I(_1387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6056__A1 (.I(_1387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6048__A1 (.I(_1387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6010__A2 (.I(_1387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8356__A1 (.I(_1390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8340__A1 (.I(_1390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8337__A1 (.I(_1390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6017__A1 (.I(_1390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6466__I (.I(_1395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6019__I (.I(_1395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6047__A2 (.I(_1397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6040__A2 (.I(_1397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6029__A2 (.I(_1397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6021__A2 (.I(_1397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8379__A1 (.I(_1400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8358__A1 (.I(_1400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7784__A1 (.I(_1400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6026__A1 (.I(_1400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6470__I (.I(_1403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6028__I (.I(_1403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7197__A2 (.I(_1404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6448__A1 (.I(_1404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6239__A2 (.I(_1404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6030__A2 (.I(_1404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8412__A1 (.I(_1406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8404__A1 (.I(_1406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7833__A1 (.I(_1406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6032__I (.I(_1406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8387__A1 (.I(_1408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8384__A1 (.I(_1408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7813__A1 (.I(_1408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6034__I (.I(_1408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8401__A1 (.I(_1409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7817__A1 (.I(_1409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7815__A1 (.I(_1409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6035__A1 (.I(_1409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6037__A2 (.I(_1410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6473__I (.I(_1413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6039__I (.I(_1413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7199__A2 (.I(_1414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6450__A1 (.I(_1414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6241__A2 (.I(_1414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6041__A2 (.I(_1414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8440__A1 (.I(_1416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8413__A1 (.I(_1416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8405__A1 (.I(_1416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6044__A1 (.I(_1416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6476__I (.I(_1419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6046__I (.I(_1419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8452__A1 (.I(_1422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8434__A1 (.I(_1422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8429__A1 (.I(_1422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6050__A1 (.I(_1422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6052__A2 (.I(_1423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8466__A1 (.I(_1429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8463__A1 (.I(_1429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8453__A1 (.I(_1429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6058__A1 (.I(_1429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6060__A2 (.I(_1430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7205__A2 (.I(_1434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6456__A1 (.I(_1434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6247__A2 (.I(_1434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6064__A2 (.I(_1434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8833__A1 (.I(_1436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8663__A1 (.I(_1436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8644__A1 (.I(_1436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6066__A1 (.I(_1436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6078__I (.I(_1437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6077__I (.I(_1437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6068__I (.I(_1437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6067__I (.I(_1437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6075__A2 (.I(_1439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6073__A2 (.I(_1439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6071__A2 (.I(_1439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6069__A2 (.I(_1439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6086__A2 (.I(_1444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6084__A2 (.I(_1444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6082__A2 (.I(_1444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6080__A2 (.I(_1444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6085__A2 (.I(_1445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6083__A2 (.I(_1445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6081__A2 (.I(_1445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6079__A2 (.I(_1445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7245__A3 (.I(_1459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6296__A2 (.I(_1459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6284__A2 (.I(_1459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6107__A1 (.I(_1459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8616__B (.I(_1460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8587__B (.I(_1460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8574__B (.I(_1460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6106__A4 (.I(_1460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8892__A2 (.I(_1461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8876__A2 (.I(_1461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6107__A2 (.I(_1461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8803__A2 (.I(_1462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6285__B (.I(_1462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6132__A1 (.I(_1462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8819__A1 (.I(_1463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7924__A2 (.I(_1463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7921__A1 (.I(_1463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6109__A1 (.I(_1463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8880__A1 (.I(_1464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6132__A2 (.I(_1464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6384__A1 (.I(_1465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6315__I (.I(_1465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6293__A1 (.I(_1465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6111__A1 (.I(_1465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8735__A1 (.I(_1466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6115__A1 (.I(_1466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6384__A2 (.I(_1467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6383__C (.I(_1467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6367__A2 (.I(_1467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6114__A1 (.I(_1467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7217__A2 (.I(_1468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6316__A2 (.I(_1468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6290__A2 (.I(_1468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6114__A2 (.I(_1468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6392__A2 (.I(_1469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6295__A3 (.I(_1469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6121__A2 (.I(_1469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6115__A2 (.I(_1469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8791__A2 (.I(_1471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6131__A1 (.I(_1471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8605__A2 (.I(_1472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8559__A2 (.I(_1472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8485__A2 (.I(_1472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6120__A2 (.I(_1472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7063__A1 (.I(_1473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6306__A1 (.I(_1473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6297__A1 (.I(_1473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6119__I (.I(_1473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8158__A1 (.I(_1474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8108__I (.I(_1474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6405__A1 (.I(_1474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6120__B (.I(_1474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8859__A2 (.I(_1476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8799__A4 (.I(_1476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6397__A2 (.I(_1476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6130__A2 (.I(_1476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8821__A1 (.I(_1477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7228__A2 (.I(_1477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6150__A1 (.I(_1477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6129__B1 (.I(_1477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8793__B (.I(_1478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6288__B (.I(_1478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6133__I (.I(_1478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6124__I (.I(_1478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8786__A1 (.I(_1479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7289__A1 (.I(_1479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6400__A1 (.I(_1479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6125__A1 (.I(_1479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7864__A1 (.I(_1481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7248__A2 (.I(_1481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7245__A2 (.I(_1481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6127__I (.I(_1481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7911__A1 (.I(_1482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7858__A3 (.I(_1482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7853__A2 (.I(_1482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6128__A4 (.I(_1482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6129__C (.I(_1483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6130__A3 (.I(_1484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6154__A2 (.I(_1487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6151__A1 (.I(_1487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8346__B2 (.I(_1488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7064__A1 (.I(_1488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6144__I (.I(_1488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6134__I (.I(_1488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8329__C (.I(_1489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8109__A1 (.I(_1489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6276__A1 (.I(_1489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6136__A1 (.I(_1489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8593__A1 (.I(_1490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7547__A1 (.I(_1490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7541__A1 (.I(_1490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6136__A2 (.I(_1490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8858__A1 (.I(_1491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6149__A2 (.I(_1491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8504__A1 (.I(_1493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8495__A1 (.I(_1493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8492__A1 (.I(_1493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6141__A1 (.I(_1493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6394__A2 (.I(_1494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6140__I (.I(_1494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8879__A2 (.I(_1495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7970__B (.I(_1495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6302__A2 (.I(_1495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6141__A2 (.I(_1495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8819__A3 (.I(_1496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6286__A2 (.I(_1496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6142__I (.I(_1496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8894__A2 (.I(_1497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8832__B2 (.I(_1497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8810__A1 (.I(_1497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6143__A2 (.I(_1497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8823__A1 (.I(_1499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7939__A2 (.I(_1499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7339__A1 (.I(_1499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6148__A1 (.I(_1499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8221__A1 (.I(_1500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7603__A2 (.I(_1500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6381__B1 (.I(_1500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6146__I (.I(_1500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8210__A1 (.I(_1501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7545__A1 (.I(_1501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6389__A2 (.I(_1501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6147__I (.I(_1501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7567__A2 (.I(_1502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7094__A1 (.I(_1502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6431__A2 (.I(_1502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6148__A2 (.I(_1502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8859__B (.I(_1503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7955__I0 (.I(_1503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6149__B2 (.I(_1503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7917__I (.I(_1507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7370__I (.I(_1507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6220__I (.I(_1507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6153__I (.I(_1507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8582__A1 (.I(_1508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6192__C (.I(_1508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6186__C (.I(_1508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6154__C (.I(_1508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8877__A2 (.I(_1509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8030__A1 (.I(_1509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7314__A2 (.I(_1509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6163__A1 (.I(_1509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8820__A1 (.I(_1510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8079__A1 (.I(_1510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8077__A1 (.I(_1510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6157__A2 (.I(_1510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8326__I (.I(_1511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8031__A2 (.I(_1511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6163__A3 (.I(_1511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8500__A2 (.I(_1512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7237__I (.I(_1512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6161__A2 (.I(_1512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7244__C (.I(_1513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6248__I (.I(_1513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6166__A1 (.I(_1513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6160__A2 (.I(_1513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7048__C (.I(_1514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6161__A4 (.I(_1514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8838__A3 (.I(_1515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6306__B (.I(_1515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6162__A3 (.I(_1515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7212__A1 (.I(_1517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6175__A1 (.I(_1517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7051__A1 (.I(_1518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7048__A1 (.I(_1518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6167__A1 (.I(_1518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7900__A3 (.I(_1519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7047__A2 (.I(_1519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6166__A2 (.I(_1519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7253__A4 (.I(_1520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7051__A2 (.I(_1520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6286__B (.I(_1520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6167__A2 (.I(_1520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6174__B (.I(_1521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6172__A1 (.I(_1521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6169__B1 (.I(_1521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6399__A2 (.I(_1524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6314__C (.I(_1524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6289__A1 (.I(_1524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6171__A1 (.I(_1524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7871__A2 (.I(_1525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6172__A2 (.I(_1525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7206__A1 (.I(_1526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6175__A3 (.I(_1526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8506__B (.I(_1528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6175__A4 (.I(_1528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6209__I (.I(_1529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6204__I (.I(_1529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6184__I (.I(_1529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6176__I (.I(_1529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8495__B (.I(_1531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7503__A2 (.I(_1531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7300__A2 (.I(_1531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6178__A2 (.I(_1531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6206__I (.I(_1532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6205__I (.I(_1532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6181__I (.I(_1532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6179__I (.I(_1532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8847__B2 (.I(_1534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8526__A1 (.I(_1534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8510__A1 (.I(_1534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6182__A1 (.I(_1534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6186__A2 (.I(_1537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8532__A1 (.I(_1540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7935__A1 (.I(_1540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7148__B2 (.I(_1540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6190__A1 (.I(_1540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8545__A1 (.I(_1541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8530__A1 (.I(_1541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8478__A1 (.I(_1541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6189__A1 (.I(_1541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6192__A2 (.I(_1543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8548__A1 (.I(_1545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7939__A1 (.I(_1545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7154__B2 (.I(_1545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6195__A1 (.I(_1545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6198__A2 (.I(_1547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8578__A1 (.I(_1550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8565__B2 (.I(_1550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8545__B2 (.I(_1550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6200__A1 (.I(_1550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6203__A2 (.I(_1552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6211__A2 (.I(_1558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8578__B2 (.I(_1561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6364__B1 (.I(_1561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6328__A1 (.I(_1561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6213__A1 (.I(_1561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6216__A2 (.I(_1563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6221__A2 (.I(_1566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7321__C (.I(_1568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7215__C (.I(_1568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6225__C (.I(_1568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6221__C (.I(_1568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6225__A2 (.I(_1570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8201__B1 (.I(_1572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8116__I (.I(_1572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8018__I (.I(_1572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6227__I (.I(_1572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8199__B1 (.I(_1573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8071__I (.I(_1573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8014__B1 (.I(_1573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6228__I (.I(_1573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8806__A2 (.I(_1574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8277__B1 (.I(_1574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8154__B1 (.I(_1574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6229__A2 (.I(_1574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6235__I (.I(_1575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6230__I (.I(_1575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6241__A1 (.I(_1577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6239__A1 (.I(_1577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6237__A1 (.I(_1577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6234__A1 (.I(_1577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6247__A1 (.I(_1578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6245__A1 (.I(_1578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6243__A1 (.I(_1578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6233__A2 (.I(_1578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6242__A2 (.I(_1580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6240__A2 (.I(_1580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6238__A2 (.I(_1580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6236__A2 (.I(_1580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7662__B (.I(_1587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7559__I (.I(_1587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7047__A1 (.I(_1587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6249__I (.I(_1587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7908__A1 (.I(_1588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7606__C (.I(_1588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7414__A1 (.I(_1588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6250__I (.I(_1588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8614__B (.I(_1589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8581__B1 (.I(_1589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8554__A1 (.I(_1589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6346__A1 (.I(_1589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6404__A1 (.I(_1590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6274__A1 (.I(_1590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6271__A1 (.I(_1590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8537__A2 (.I(_1591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6253__A2 (.I(_1591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6274__A3 (.I(_1594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6263__A2 (.I(_1601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6268__A2 (.I(_1602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6273__A2 (.I(_1611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8847__C (.I(_1614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8836__A1 (.I(_1614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6406__A1 (.I(_1614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6276__A2 (.I(_1614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8619__B1 (.I(_1615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8530__A2 (.I(_1615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8510__A2 (.I(_1615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6345__A1 (.I(_1615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6279__A1 (.I(_1616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6279__A2 (.I(_1617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6314__A2 (.I(_1618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6282__A2 (.I(_1618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8607__B2 (.I(_1619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6407__A1 (.I(_1619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6330__A1 (.I(_1619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6281__A1 (.I(_1619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8879__A1 (.I(_1622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8416__B (.I(_1622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6295__A2 (.I(_1622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6286__A1 (.I(_1622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8867__A1 (.I(_1626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8842__B (.I(_1626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7855__A1 (.I(_1626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6289__A2 (.I(_1626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8508__A1 (.I(_1628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6308__A1 (.I(_1628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7226__A3 (.I(_1629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6291__B (.I(_1629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8844__A1 (.I(_1630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8801__A1 (.I(_1630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8502__B (.I(_1630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6292__B (.I(_1630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8868__A2 (.I(_1631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6308__A2 (.I(_1631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8703__A1 (.I(_1633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7002__A1 (.I(_1633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7000__A1 (.I(_1633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6295__A1 (.I(_1633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8839__A3 (.I(_1634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6298__A1 (.I(_1634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8501__C (.I(_1635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7224__A1 (.I(_1635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6298__A2 (.I(_1635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8841__C (.I(_1636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6298__A3 (.I(_1636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8526__C (.I(_1639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6402__B (.I(_1639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6357__I (.I(_1639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6301__A2 (.I(_1639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8591__A1 (.I(_1640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8539__I (.I(_1640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6302__A4 (.I(_1640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8507__A1 (.I(_1642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6307__B1 (.I(_1642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8805__I (.I(_1643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8501__A2 (.I(_1643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7251__A1 (.I(_1643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6305__A1 (.I(_1643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8832__A1 (.I(_1644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8830__A2 (.I(_1644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6306__A2 (.I(_1644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6307__C (.I(_1645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6409__S (.I(_1648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6349__A2 (.I(_1648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6345__B (.I(_1648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7249__A1 (.I(_1649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6311__I (.I(_1649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8578__A2 (.I(_1650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6326__A2 (.I(_1650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6325__A1 (.I(_1650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6312__A1 (.I(_1650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8892__A1 (.I(_1654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7970__C (.I(_1654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6383__A1 (.I(_1654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6324__A1 (.I(_1654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8237__A1 (.I(_1657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7791__A2 (.I(_1657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7579__A1 (.I(_1657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6319__I (.I(_1657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6389__B1 (.I(_1658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6377__B1 (.I(_1658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6322__A2 (.I(_1658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6320__I (.I(_1658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8608__A1 (.I(_1659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7097__A1 (.I(_1659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6929__A1 (.I(_1659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6323__A2 (.I(_1659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8603__A1 (.I(_1660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6377__B2 (.I(_1660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6349__A1 (.I(_1660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6322__A1 (.I(_1660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6324__A4 (.I(_1662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6326__C (.I(_1664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8589__B2 (.I(_1668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6903__A1 (.I(_1668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6361__A1 (.I(_1668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6330__A4 (.I(_1668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6332__A3 (.I(_1669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8172__A1 (.I(_1672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7514__A2 (.I(_1672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7087__I (.I(_1672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6336__A1 (.I(_1672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7611__A2 (.I(_1673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7592__A1 (.I(_1673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7584__A1 (.I(_1673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6335__I (.I(_1673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8244__A1 (.I(_1674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7959__A2 (.I(_1674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6434__A1 (.I(_1674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6336__A3 (.I(_1674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8004__A1 (.I(_1676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7928__A2 (.I(_1676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6415__I (.I(_1676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6342__A1 (.I(_1676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8823__A2 (.I(_1677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8527__A1 (.I(_1677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6424__A2 (.I(_1677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6342__A2 (.I(_1677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8546__A1 (.I(_1678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7940__A2 (.I(_1678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6427__A1 (.I(_1678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6342__A3 (.I(_1678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8143__A1 (.I(_1679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7434__A1 (.I(_1679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6368__A1 (.I(_1679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6341__I (.I(_1679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8781__A1 (.I(_1680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8137__A1 (.I(_1680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7944__A2 (.I(_1680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6342__A4 (.I(_1680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6344__B1 (.I(_1682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6345__C (.I(_1683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6350__A1 (.I(_1685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8123__I (.I(_1686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7220__I (.I(_1686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6351__I (.I(_1686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6348__I (.I(_1686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8083__A1 (.I(_1687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8037__B (.I(_1687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7529__B (.I(_1687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6349__B (.I(_1687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8826__A1 (.I(_1689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7419__A1 (.I(_1689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7231__C (.I(_1689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6410__A1 (.I(_1689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8615__A1 (.I(_1690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6409__I0 (.I(_1690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6398__B2 (.I(_1690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6395__A1 (.I(_1690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8871__A1 (.I(_1691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8529__A1 (.I(_1691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8490__B (.I(_1691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6408__A1 (.I(_1691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8250__A1 (.I(_1692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8094__A2 (.I(_1692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6397__A1 (.I(_1692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6355__I (.I(_1692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8362__A1 (.I(_1693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8026__A1 (.I(_1693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7521__A1 (.I(_1693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6356__I (.I(_1693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7970__A2 (.I(_1694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7776__A1 (.I(_1694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7404__A1 (.I(_1694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6403__A1 (.I(_1694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8527__A2 (.I(_1695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8489__A2 (.I(_1695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8488__A1 (.I(_1695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6403__A2 (.I(_1695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8618__B (.I(_1699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6402__A1 (.I(_1699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8588__C (.I(_1700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8543__B (.I(_1700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8486__C (.I(_1700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6363__I (.I(_1700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8576__B (.I(_1701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8555__I (.I(_1701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8525__B (.I(_1701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6401__A1 (.I(_1701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6383__B (.I(_1704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6367__A3 (.I(_1704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6368__C (.I(_1705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6393__A1 (.I(_1707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7309__A1 (.I(_1708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7035__I (.I(_1708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6386__A2 (.I(_1708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6373__B1 (.I(_1708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7445__A2 (.I(_1709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6386__B1 (.I(_1709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6372__I (.I(_1709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7467__A2 (.I(_1710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7423__A1 (.I(_1710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7083__I (.I(_1710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6373__C2 (.I(_1710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6382__A1 (.I(_1711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7356__A1 (.I(_1712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6387__A2 (.I(_1712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6375__I (.I(_1712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7359__A1 (.I(_1713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7354__A1 (.I(_1713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7073__I (.I(_1713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6377__A2 (.I(_1713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7447__A2 (.I(_1717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7424__A1 (.I(_1717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7384__B (.I(_1717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6380__I (.I(_1717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7393__A1 (.I(_1718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7078__I (.I(_1718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6387__B1 (.I(_1718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6381__A2 (.I(_1718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6383__A2 (.I(_1720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6389__C (.I(_1726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6390__A4 (.I(_1727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8734__A1 (.I(_1729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6538__A1 (.I(_1729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6513__A1 (.I(_1729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6392__A1 (.I(_1729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6395__A3 (.I(_1730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6393__C (.I(_1730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6398__A1 (.I(_1731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8882__A1 (.I(_1732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8870__A1 (.I(_1732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8846__A1 (.I(_1732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6396__A1 (.I(_1732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7963__A1 (.I(_1737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6406__A2 (.I(_1737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6400__B (.I(_1737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6408__A2 (.I(_1741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6408__B1 (.I(_1742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6408__B2 (.I(_1745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6409__I1 (.I(_1746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7902__A2 (.I(_1749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7252__B (.I(_1749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6413__A2 (.I(_1749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6436__A2 (.I(_1751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6434__A2 (.I(_1751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6427__A2 (.I(_1751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6423__A1 (.I(_1751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8828__A2 (.I(_1752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8489__A1 (.I(_1752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7303__A1 (.I(_1752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6416__A2 (.I(_1752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8783__A2 (.I(_1754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8781__A2 (.I(_1754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6425__I (.I(_1754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6421__A1 (.I(_1754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8463__A2 (.I(_1755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6419__A2 (.I(_1755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8794__B1 (.I(_1756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8455__B (.I(_1756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6420__A4 (.I(_1756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6421__A2 (.I(_1757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6436__B1 (.I(_1758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6434__B1 (.I(_1758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6422__I (.I(_1758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8784__A2 (.I(_1761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8782__A2 (.I(_1761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6433__A2 (.I(_1761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6426__B2 (.I(_1761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6428__I (.I(_1762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8497__A1 (.I(_1764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7412__A1 (.I(_1764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7040__A2 (.I(_1764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6432__A2 (.I(_1764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6432__B (.I(_1765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6433__B2 (.I(_1766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6437__I (.I(_1768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6444__I (.I(_1769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6439__I (.I(_1769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6455__A2 (.I(_1770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6453__A2 (.I(_1770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6441__I (.I(_1770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6440__I (.I(_1770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6450__A2 (.I(_1771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6448__A2 (.I(_1771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6446__A2 (.I(_1771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6443__A2 (.I(_1771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6456__A2 (.I(_1772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6454__A2 (.I(_1772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6452__A2 (.I(_1772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6442__A2 (.I(_1772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6451__A2 (.I(_1774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6449__A2 (.I(_1774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6447__A2 (.I(_1774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6445__A2 (.I(_1774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8689__A1 (.I(_1781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8649__A1 (.I(_1781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7110__A1 (.I(_1781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6465__A1 (.I(_1781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8684__A3 (.I(_1782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8644__A2 (.I(_1782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7105__A3 (.I(_1782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6460__A2 (.I(_1782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6467__I (.I(_1784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6461__I (.I(_1784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6483__A2 (.I(_1785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6480__A2 (.I(_1785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6463__I (.I(_1785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6462__I (.I(_1785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6475__A2 (.I(_1786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6472__A2 (.I(_1786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6469__A2 (.I(_1786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6465__A2 (.I(_1786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6484__A2 (.I(_1787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6481__A2 (.I(_1787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6478__A2 (.I(_1787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6464__A2 (.I(_1787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8692__A1 (.I(_1789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8652__A1 (.I(_1789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7113__A1 (.I(_1789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6469__A1 (.I(_1789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6477__A2 (.I(_1790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6474__A2 (.I(_1790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6471__A2 (.I(_1790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6468__A2 (.I(_1790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8694__A1 (.I(_1792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8654__A1 (.I(_1792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7115__A1 (.I(_1792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6472__A1 (.I(_1792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8696__A1 (.I(_1794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8656__A1 (.I(_1794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7117__A1 (.I(_1794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6475__A1 (.I(_1794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8698__A1 (.I(_1796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8658__A1 (.I(_1796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7119__A1 (.I(_1796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6478__A1 (.I(_1796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8700__A1 (.I(_1798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8660__A1 (.I(_1798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7121__A1 (.I(_1798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6481__A1 (.I(_1798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8702__A1 (.I(_1800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8662__A1 (.I(_1800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7123__A1 (.I(_1800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6484__A1 (.I(_1800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7922__A1 (.I(_1802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6488__A2 (.I(_1802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6507__A3 (.I(_1803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6487__I (.I(_1803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6518__I (.I(_1805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6489__I (.I(_1805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6783__I (.I(_1806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6727__I (.I(_1806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6530__A1 (.I(_1806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6511__B (.I(_1806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7130__A3 (.I(_1808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6523__A2 (.I(_1808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6502__A2 (.I(_1808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6492__A3 (.I(_1808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6955__C (.I(_1810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6524__B (.I(_1810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6494__I (.I(_1810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6899__A2 (.I(_1812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6743__A2 (.I(_1812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6536__A2 (.I(_1812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6496__A2 (.I(_1812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6831__A2 (.I(_1813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6733__I (.I(_1813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6520__I (.I(_1813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6497__I (.I(_1813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6929__A2 (.I(_1814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6888__A2 (.I(_1814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6788__A2 (.I(_1814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6510__A2 (.I(_1814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7136__A2 (.I(_1815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7133__A2 (.I(_1815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7126__A2 (.I(_1815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6499__A2 (.I(_1815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6956__B (.I(_1817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6785__I (.I(_1817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6729__I (.I(_1817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6501__I (.I(_1817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6903__B (.I(_1818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6833__B (.I(_1818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6736__B (.I(_1818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6505__A1 (.I(_1818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6533__I (.I(_1819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6505__A2 (.I(_1819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6519__I (.I(_1820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6504__I (.I(_1820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6516__I (.I(_1825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6509__I (.I(_1825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6908__A2 (.I(_1826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6894__A2 (.I(_1826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6794__A2 (.I(_1826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6510__A4 (.I(_1826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6511__C (.I(_1827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7125__A2 (.I(_1828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6512__I (.I(_1828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6897__A1 (.I(_1830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6514__I (.I(_1830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6969__A1 (.I(_1831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6952__A1 (.I(_1831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6926__A1 (.I(_1831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6515__I (.I(_1831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6865__A1 (.I(_1832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6829__A1 (.I(_1832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6780__A1 (.I(_1832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6723__A1 (.I(_1832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6782__I (.I(_1833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6724__I (.I(_1833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6531__B (.I(_1833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6517__I (.I(_1833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6905__B (.I(_1835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6791__B (.I(_1835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6725__I (.I(_1835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6531__A2 (.I(_1835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6957__C (.I(_1836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6834__B (.I(_1836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6726__I (.I(_1836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6529__A2 (.I(_1836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8490__A2 (.I(_1839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6524__A1 (.I(_1839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6955__A2 (.I(_1840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6954__A2 (.I(_1840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6928__A2 (.I(_1840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6524__A2 (.I(_1840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6932__A1 (.I(_1842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6931__A2 (.I(_1842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6527__A2 (.I(_1842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6526__C (.I(_1842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6961__C (.I(_1850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6781__I (.I(_1850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6741__I (.I(_1850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6534__S (.I(_1850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6535__I (.I(_1851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7139__A1 (.I(_1852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7005__A1 (.I(_1852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6723__A2 (.I(_1852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7144__I (.I(_1853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6720__I (.I(_1853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6537__I (.I(_1853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7137__A1 (.I(_1854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7025__I (.I(_1854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7002__B (.I(_1854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6538__B (.I(_1854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6968__A2 (.I(_1856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6898__A2 (.I(_1856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6779__A2 (.I(_1856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6722__A2 (.I(_1856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6767__A2 (.I(_1857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6710__A2 (.I(_1857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6631__A2 (.I(_1857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6541__I (.I(_1857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6769__A2 (.I(_1860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6671__A2 (.I(_1860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6632__A2 (.I(_1860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6544__I (.I(_1860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6662__A1 (.I(_1863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6660__A1 (.I(_1863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6630__A1 (.I(_1863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6550__A1 (.I(_1863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8588__A1 (.I(_1864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6870__A2 (.I(_1864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6844__A2 (.I(_1864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6549__A2 (.I(_1864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8576__A1 (.I(_1865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6846__A2 (.I(_1865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6562__A2 (.I(_1865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6549__B1 (.I(_1865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6636__A2 (.I(_1868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6552__I (.I(_1868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6578__I (.I(_1871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6555__I (.I(_1871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6697__A1 (.I(_1873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6626__A1 (.I(_1873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6560__A2 (.I(_1873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6653__A2 (.I(_1874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6635__A2 (.I(_1874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6625__A2 (.I(_1874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6558__I (.I(_1874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6626__A2 (.I(_1876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6584__A1 (.I(_1876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6560__A3 (.I(_1876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6623__A1 (.I(_1878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6622__A1 (.I(_1878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6576__A1 (.I(_1878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6654__A1 (.I(_1881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6570__A1 (.I(_1881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6569__A1 (.I(_1881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6567__A2 (.I(_1881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6704__A2 (.I(_1882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6598__I (.I(_1882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6583__A2 (.I(_1882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6566__A2 (.I(_1882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6650__A2 (.I(_1889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6573__I (.I(_1889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6621__A2 (.I(_1891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6575__A2 (.I(_1891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6703__A2 (.I(_1895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6637__A2 (.I(_1895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6597__A2 (.I(_1895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6579__I (.I(_1895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6605__I (.I(_1896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6593__A3 (.I(_1896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6583__B1 (.I(_1896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6580__A2 (.I(_1896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7008__A1 (.I(_1897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6584__A2 (.I(_1897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6610__A4 (.I(_1898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6606__I (.I(_1898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6593__A4 (.I(_1898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6582__A2 (.I(_1898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6758__A2 (.I(_1902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6594__A2 (.I(_1902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6588__I (.I(_1902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6586__A2 (.I(_1902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6688__I (.I(_1906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6647__A2 (.I(_1906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6608__A2 (.I(_1906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6590__A2 (.I(_1906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8559__A1 (.I(_1915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6851__A2 (.I(_1915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6808__A2 (.I(_1915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6599__A2 (.I(_1915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8524__A1 (.I(_1922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6612__A2 (.I(_1922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6610__A3 (.I(_1922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6608__A3 (.I(_1922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8485__A1 (.I(_1923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7007__A2 (.I(_1923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6612__B1 (.I(_1923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6607__A2 (.I(_1923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8709__A2 (.I(_1924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7004__A2 (.I(_1924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6608__A4 (.I(_1924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7028__A2 (.I(_1937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7024__A1 (.I(_1937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6644__A2 (.I(_1937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6696__A1 (.I(_1942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6666__A1 (.I(_1942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6627__A1 (.I(_1942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6649__A1 (.I(_1946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6641__A1 (.I(_1946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6648__A2 (.I(_1956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6640__A2 (.I(_1956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6684__A1 (.I(_1964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6678__A1 (.I(_1964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6815__A1 (.I(_1968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6769__A1 (.I(_1968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6653__B2 (.I(_1968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6652__A1 (.I(_1968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6756__A2 (.I(_1973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6698__A2 (.I(_1973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6686__I (.I(_1973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6657__A2 (.I(_1973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6702__A1 (.I(_1983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6675__A1 (.I(_1983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6692__A2 (.I(_1992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6691__A2 (.I(_1992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6676__A3 (.I(_1992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6842__I (.I(_2003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6807__A2 (.I(_2003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6750__A2 (.I(_2003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6687__A2 (.I(_2003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8542__A1 (.I(_2005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6802__A2 (.I(_2005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6751__A2 (.I(_2005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6689__A2 (.I(_2005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6755__A1 (.I(_2017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6715__A1 (.I(_2017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6820__A1 (.I(_2021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6803__A2 (.I(_2021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6705__A2 (.I(_2021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6761__A2 (.I(_2030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6714__A2 (.I(_2030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6746__A2 (.I(_2034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6718__A2 (.I(_2034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8738__A2 (.I(_2036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6722__B1 (.I(_2036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7170__A1 (.I(_2037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7010__I (.I(_2037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6827__I (.I(_2037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6721__I (.I(_2037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7004__A1 (.I(_2038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6967__A1 (.I(_2038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6779__B2 (.I(_2038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6722__B2 (.I(_2038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6787__I (.I(_2046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6731__I (.I(_2046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6909__A2 (.I(_2059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6908__B (.I(_2059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6886__A2 (.I(_2059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6744__A2 (.I(_2059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7149__A1 (.I(_2061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7012__A1 (.I(_2061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6780__A2 (.I(_2061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6798__A1 (.I(_2065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6777__A1 (.I(_2065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6762__A1 (.I(_2076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6808__A3 (.I(_2087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6772__A2 (.I(_2087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6798__A2 (.I(_2092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6777__A2 (.I(_2092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6960__A2 (.I(_2098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6906__A2 (.I(_2098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6892__A1 (.I(_2098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6792__A2 (.I(_2098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7155__A1 (.I(_2111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7015__A1 (.I(_2111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6829__A2 (.I(_2111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6951__A2 (.I(_2112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6925__A2 (.I(_2112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6864__A2 (.I(_2112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6828__A2 (.I(_2112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6861__A1 (.I(_2116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6825__A1 (.I(_2116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6841__A1 (.I(_2118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6824__A1 (.I(_2118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6840__A1 (.I(_2121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6823__A1 (.I(_2121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6840__A2 (.I(_2137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6823__A2 (.I(_2137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8746__A2 (.I(_2141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6828__B1 (.I(_2141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6951__B2 (.I(_2142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6925__B2 (.I(_2142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6864__B2 (.I(_2142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6828__B2 (.I(_2142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8589__A1 (.I(_2144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8581__A1 (.I(_2144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8563__B2 (.I(_2144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6833__A1 (.I(_2144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7160__A1 (.I(_2153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7018__A1 (.I(_2153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6865__A2 (.I(_2153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6866__A1 (.I(_2168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6857__A1 (.I(_2168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6866__A2 (.I(_2170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6857__A2 (.I(_2170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6883__B (.I(_2172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6860__A1 (.I(_2172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8748__A2 (.I(_2177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6864__B1 (.I(_2177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6921__B2 (.I(_2180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6877__A1 (.I(_2180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6911__A1 (.I(_2190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6881__A1 (.I(_2190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6911__A2 (.I(_2193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6881__A2 (.I(_2193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8751__A3 (.I(_2198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6899__A3 (.I(_2198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6896__A2 (.I(_2208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7166__A1 (.I(_2209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7022__A1 (.I(_2209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6897__A2 (.I(_2209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6910__I (.I(_2221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7171__A1 (.I(_2222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7027__A1 (.I(_2222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6926__A2 (.I(_2222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8617__A1 (.I(_2230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6945__A2 (.I(_2230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6944__A2 (.I(_2230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6919__A2 (.I(_2230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6938__A2 (.I(_2235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6937__A2 (.I(_2235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6924__A3 (.I(_2235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7177__A1 (.I(_2247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7031__A1 (.I(_2247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6952__A2 (.I(_2247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6966__A2 (.I(_2260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6950__A2 (.I(_2260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8755__A2 (.I(_2261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6951__B1 (.I(_2261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8141__A1 (.I(_2263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8057__A1 (.I(_2263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7669__A1 (.I(_2263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6954__A1 (.I(_2263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7181__A1 (.I(_2272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7034__A1 (.I(_2272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6969__A2 (.I(_2272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6966__B (.I(_2275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8758__A2 (.I(_2276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6967__A2 (.I(_2276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8764__A1 (.I(_2279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8667__A1 (.I(_2279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8627__A1 (.I(_2279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6976__A1 (.I(_2279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8813__A1 (.I(_2280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8760__A1 (.I(_2280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8663__A3 (.I(_2280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6972__A1 (.I(_2280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6988__I (.I(_2281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6987__I (.I(_2281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6974__I (.I(_2281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6973__I (.I(_2281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6984__A2 (.I(_2283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6981__A2 (.I(_2283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6978__A2 (.I(_2283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6975__A2 (.I(_2283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8766__A1 (.I(_2285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8669__A1 (.I(_2285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8629__A1 (.I(_2285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6979__A1 (.I(_2285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8768__A1 (.I(_2287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8671__A1 (.I(_2287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8631__A1 (.I(_2287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6982__A1 (.I(_2287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8770__A1 (.I(_2289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8673__A1 (.I(_2289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8633__A1 (.I(_2289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6985__A1 (.I(_2289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8774__A1 (.I(_2291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8677__A1 (.I(_2291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8637__A1 (.I(_2291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6990__A1 (.I(_2291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8776__A1 (.I(_2295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8679__A1 (.I(_2295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8639__A1 (.I(_2295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6993__A1 (.I(_2295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8778__A1 (.I(_2297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8681__A1 (.I(_2297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8641__A1 (.I(_2297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6996__A1 (.I(_2297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8780__A1 (.I(_2299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8683__A1 (.I(_2299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8643__A1 (.I(_2299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6999__A1 (.I(_2299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7018__A2 (.I(_2302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7015__A2 (.I(_2302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7012__A2 (.I(_2302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7005__A2 (.I(_2302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7006__I (.I(_2303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7003__I (.I(_2303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7033__A2 (.I(_2304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7030__A2 (.I(_2304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7026__A2 (.I(_2304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7004__B1 (.I(_2304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8715__A2 (.I(_2309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7011__B1 (.I(_2309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8718__A2 (.I(_2312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7014__B1 (.I(_2312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8720__A2 (.I(_2314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7017__B1 (.I(_2314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7034__A2 (.I(_2316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7031__A2 (.I(_2316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7027__A2 (.I(_2316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7022__A2 (.I(_2316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8723__A2 (.I(_2317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7021__B1 (.I(_2317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8727__A2 (.I(_2320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7026__B1 (.I(_2320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7176__A1 (.I(_2321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7033__B2 (.I(_2321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7030__B2 (.I(_2321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7026__B2 (.I(_2321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8730__A2 (.I(_2324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7030__B1 (.I(_2324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8732__A2 (.I(_2326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7033__B1 (.I(_2326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7312__B (.I(_2328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7296__A2 (.I(_2328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7279__A2 (.I(_2328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7036__I (.I(_2328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8319__A1 (.I(_2329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7997__B2 (.I(_2329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7307__A1 (.I(_2329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7072__A1 (.I(_2329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8211__B2 (.I(_2330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8049__B2 (.I(_2330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7738__I (.I(_2330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7038__I (.I(_2330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8006__A2 (.I(_2331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7781__B1 (.I(_2331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7641__C (.I(_2331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7040__A1 (.I(_2331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7260__A2 (.I(_2332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7040__A3 (.I(_2332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8209__A2 (.I(_2334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8055__A2 (.I(_2334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7894__A2 (.I(_2334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7042__I (.I(_2334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8172__A2 (.I(_2335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7779__B (.I(_2335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7408__I (.I(_2335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7044__A2 (.I(_2335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8790__B (.I(_2336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8787__A2 (.I(_2336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7782__I (.I(_2336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7044__A3 (.I(_2336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7243__B1 (.I(_2338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7046__A2 (.I(_2338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8497__B (.I(_2341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7058__A1 (.I(_2341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7881__A3 (.I(_2342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7057__A1 (.I(_2342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8837__A2 (.I(_2343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8502__A2 (.I(_2343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7206__A2 (.I(_2343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7057__A2 (.I(_2343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8506__A1 (.I(_2344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8494__A2 (.I(_2344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7858__A4 (.I(_2344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7055__A1 (.I(_2344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7436__I (.I(_2345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7353__I (.I(_2345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7053__A2 (.I(_2345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7553__I (.I(_2346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7361__I (.I(_2346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7054__A2 (.I(_2346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7400__A1 (.I(_2347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7316__A2 (.I(_2347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7055__A2 (.I(_2347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7057__A3 (.I(_2348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7065__A3 (.I(_2351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8500__A1 (.I(_2352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8001__A1 (.I(_2352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7882__I (.I(_2352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7060__A1 (.I(_2352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8368__B (.I(_2354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8173__C (.I(_2354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8138__C (.I(_2354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7064__B1 (.I(_2354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8363__A2 (.I(_2355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8236__I (.I(_2355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7410__B (.I(_2355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7063__A2 (.I(_2355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7100__A2 (.I(_2359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7096__A2 (.I(_2359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7090__S (.I(_2359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7067__I (.I(_2359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7086__A2 (.I(_2360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7082__A2 (.I(_2360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7077__A2 (.I(_2360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7072__A2 (.I(_2360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8318__A1 (.I(_2361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7676__A1 (.I(_2361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7671__A1 (.I(_2361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7069__I (.I(_2361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8317__A1 (.I(_2362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7998__A1 (.I(_2362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7694__A2 (.I(_2362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7071__A1 (.I(_2362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7101__A2 (.I(_2363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7097__A2 (.I(_2363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7094__A2 (.I(_2363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7071__A2 (.I(_2363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8819__A2 (.I(_2365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7936__A2 (.I(_2365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7343__A2 (.I(_2365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7077__A1 (.I(_2365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8366__A2 (.I(_2366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8343__A1 (.I(_2366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8063__B2 (.I(_2366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7076__A1 (.I(_2366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7093__A2 (.I(_2367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7085__A2 (.I(_2367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7081__A2 (.I(_2367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7076__A2 (.I(_2367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8364__A1 (.I(_2369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8098__A1 (.I(_2369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8093__A1 (.I(_2369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7082__A1 (.I(_2369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8367__A1 (.I(_2370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8363__A1 (.I(_2370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7778__A2 (.I(_2370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7080__I (.I(_2370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8368__A1 (.I(_2371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7757__A1 (.I(_2371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7754__A1 (.I(_2371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7081__A1 (.I(_2371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8565__A1 (.I(_2373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7437__A1 (.I(_2373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7430__A1 (.I(_2373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7086__A1 (.I(_2373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8437__A1 (.I(_2374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8393__A1 (.I(_2374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8388__A1 (.I(_2374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7085__A1 (.I(_2374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8579__A1 (.I(_2376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7505__A1 (.I(_2376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7496__A1 (.I(_2376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7088__I (.I(_2376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8875__A2 (.I(_2377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8783__A1 (.I(_2377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7950__A2 (.I(_2377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7090__I0 (.I(_2377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8437__A2 (.I(_2378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8410__A1 (.I(_2378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8408__A1 (.I(_2378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7090__I1 (.I(_2378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8436__A1 (.I(_2380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8435__A1 (.I(_2380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7912__A1 (.I(_2380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7093__A1 (.I(_2380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8460__A1 (.I(_2382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8252__B2 (.I(_2382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7915__A1 (.I(_2382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7096__A1 (.I(_2382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8414__A1 (.I(_2384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7639__A2 (.I(_2384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7282__I (.I(_2384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7099__I (.I(_2384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8619__A1 (.I(_2385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8329__A1 (.I(_2385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7898__A1 (.I(_2385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7101__A1 (.I(_2385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8017__I (.I(_2387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8013__I (.I(_2387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7103__I (.I(_2387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8184__A2 (.I(_2388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8182__A2 (.I(_2388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8117__A2 (.I(_2388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7104__I (.I(_2388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8281__A2 (.I(_2389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8277__A2 (.I(_2389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8153__A2 (.I(_2389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7105__A2 (.I(_2389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7122__A2 (.I(_2391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7120__A2 (.I(_2391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7108__I (.I(_2391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7107__I (.I(_2391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7117__A2 (.I(_2392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7115__A2 (.I(_2392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7113__A2 (.I(_2392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7110__A2 (.I(_2392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7123__A2 (.I(_2393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7121__A2 (.I(_2393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7119__A2 (.I(_2393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7109__A2 (.I(_2393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7118__A2 (.I(_2395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7116__A2 (.I(_2395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7114__A2 (.I(_2395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7112__A2 (.I(_2395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8605__B1 (.I(_2402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8558__B (.I(_2402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7136__A1 (.I(_2402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7126__A1 (.I(_2402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7142__I (.I(_2403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7128__I (.I(_2403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7126__B (.I(_2403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8225__A1 (.I(_2407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7957__I (.I(_2407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7933__I (.I(_2407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7130__A1 (.I(_2407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7152__I (.I(_2408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7131__I (.I(_2408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7180__A2 (.I(_2409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7175__A2 (.I(_2409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7147__A2 (.I(_2409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7135__A2 (.I(_2409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8818__A1 (.I(_2410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8575__A1 (.I(_2410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8520__A1 (.I(_2410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7133__A1 (.I(_2410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7165__A1 (.I(_2421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7159__A1 (.I(_2421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7154__A1 (.I(_2421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7148__A1 (.I(_2421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7165__C (.I(_2438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8008__I (.I(_2454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7185__I (.I(_2454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8200__A2 (.I(_2455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8185__A2 (.I(_2455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8151__A2 (.I(_2455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7186__I (.I(_2455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8278__A2 (.I(_2456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8155__A2 (.I(_2456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8073__A2 (.I(_2456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7187__A2 (.I(_2456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7193__I (.I(_2457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7188__I (.I(_2457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7204__A2 (.I(_2458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7202__A2 (.I(_2458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7190__I (.I(_2458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7189__I (.I(_2458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7199__A1 (.I(_2459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7197__A1 (.I(_2459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7195__A1 (.I(_2459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7192__A1 (.I(_2459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7205__A1 (.I(_2460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7203__A1 (.I(_2460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7201__A1 (.I(_2460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7191__A2 (.I(_2460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7200__A2 (.I(_2462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7198__A2 (.I(_2462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7196__A2 (.I(_2462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7194__A2 (.I(_2462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8790__A1 (.I(_2471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8027__I (.I(_2471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7285__A1 (.I(_2471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7209__I (.I(_2471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8842__A2 (.I(_2472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8444__A1 (.I(_2472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8157__A1 (.I(_2472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7210__I (.I(_2472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8828__A1 (.I(_2473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8421__A1 (.I(_2473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7932__I (.I(_2473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7211__A1 (.I(_2473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7215__A1 (.I(_2475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7214__A2 (.I(_2475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7215__A2 (.I(_2476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7915__A2 (.I(_2478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7912__A2 (.I(_2478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7268__A2 (.I(_2478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7218__A1 (.I(_2478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7224__A2 (.I(_2479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7218__A2 (.I(_2479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7978__C (.I(_2480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7262__A1 (.I(_2480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7219__A3 (.I(_2480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7222__A2 (.I(_2481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7221__A2 (.I(_2481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8596__B (.I(_2482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8532__B (.I(_2482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8514__B (.I(_2482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7221__B (.I(_2482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7901__C (.I(_2486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7888__A3 (.I(_2486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7860__A4 (.I(_2486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7226__A2 (.I(_2486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7885__A2 (.I(_2487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7859__A1 (.I(_2487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7229__A3 (.I(_2487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7980__B1 (.I(_2488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7228__A4 (.I(_2488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7861__A1 (.I(_2489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7229__A4 (.I(_2489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7883__A2 (.I(_2494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7856__A3 (.I(_2494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7252__A2 (.I(_2494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7235__A2 (.I(_2494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7866__A2 (.I(_2496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7263__A1 (.I(_2496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8376__A1 (.I(_2497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8260__I (.I(_2497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7981__A1 (.I(_2497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7239__A1 (.I(_2497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8877__A3 (.I(_2498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7975__A2 (.I(_2498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7881__A1 (.I(_2498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7239__A2 (.I(_2498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7861__A2 (.I(_2499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7263__A2 (.I(_2499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7892__A1 (.I(_2500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7263__A3 (.I(_2500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7243__B2 (.I(_2502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7891__A1 (.I(_2503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7247__A1 (.I(_2503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7910__A1 (.I(_2504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7247__A2 (.I(_2504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7247__A3 (.I(_2505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7973__I (.I(_2510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7972__C (.I(_2510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7251__C (.I(_2510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7854__A1 (.I(_2511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7261__A1 (.I(_2511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7910__A2 (.I(_2512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7862__I (.I(_2512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7254__A1 (.I(_2512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7910__A3 (.I(_2513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7254__A2 (.I(_2513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7256__A2 (.I(_2515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7257__B (.I(_2516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7854__A2 (.I(_2517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7261__A3 (.I(_2517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7878__A3 (.I(_2518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7875__A3 (.I(_2518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7874__A2 (.I(_2518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7259__A2 (.I(_2518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7263__A4 (.I(_2522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7417__I (.I(_2523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7264__I (.I(_2523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7574__I (.I(_2524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7531__I (.I(_2524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7322__I (.I(_2524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7265__I (.I(_2524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7852__A1 (.I(_2526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7819__A1 (.I(_2526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7790__A1 (.I(_2526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7321__A1 (.I(_2526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8037__A1 (.I(_2527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8033__A1 (.I(_2527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7319__A1 (.I(_2527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7275__A1 (.I(_2527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7561__I (.I(_2528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7525__I (.I(_2528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7474__I (.I(_2528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7269__A2 (.I(_2528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7627__I (.I(_2529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7475__A2 (.I(_2529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7324__I (.I(_2529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7270__I (.I(_2529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7850__A2 (.I(_2530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7817__A2 (.I(_2530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7573__A2 (.I(_2530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7319__A2 (.I(_2530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8322__A1 (.I(_2531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8253__A1 (.I(_2531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7846__A2 (.I(_2531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7273__A1 (.I(_2531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7619__A2 (.I(_2533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7473__A2 (.I(_2533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7407__A3 (.I(_2533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7274__I (.I(_2533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7708__A2 (.I(_2534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7571__A2 (.I(_2534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7524__A2 (.I(_2534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7318__A1 (.I(_2534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8384__A2 (.I(_2538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8328__A2 (.I(_2538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7334__A2 (.I(_2538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7287__A1 (.I(_2538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8026__A2 (.I(_2539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7996__A2 (.I(_2539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7315__A2 (.I(_2539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7287__A2 (.I(_2539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7320__A1 (.I(_2541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7316__A1 (.I(_2541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7298__A1 (.I(_2541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7283__A1 (.I(_2541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7842__A2 (.I(_2542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7809__A2 (.I(_2542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7735__A2 (.I(_2542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7283__A2 (.I(_2542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7775__B (.I(_2546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7403__B (.I(_2546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7335__A1 (.I(_2546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7287__C (.I(_2546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8350__C (.I(_2548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8224__C (.I(_2548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8188__B (.I(_2548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7289__A3 (.I(_2548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7345__C (.I(_2549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7298__B (.I(_2549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7810__A1 (.I(_2550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7736__A1 (.I(_2550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7639__A1 (.I(_2550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7291__I (.I(_2550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7694__A1 (.I(_2551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7409__A1 (.I(_2551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7344__A2 (.I(_2551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7297__A2 (.I(_2551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8296__A1 (.I(_2552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8222__A2 (.I(_2552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7341__I (.I(_2552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7293__I (.I(_2552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8388__A2 (.I(_2553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7812__A1 (.I(_2553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7739__A1 (.I(_2553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7297__B (.I(_2553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8290__A1 (.I(_2554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7566__I (.I(_2554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7342__I (.I(_2554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7295__I (.I(_2554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7858__A1 (.I(_2555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7778__A1 (.I(_2555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7514__A1 (.I(_2555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7296__A1 (.I(_2555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7297__C (.I(_2556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7352__A1 (.I(_2560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7304__I (.I(_2560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7301__I (.I(_2560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7657__A1 (.I(_2562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7546__A1 (.I(_2562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7502__A1 (.I(_2562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7303__A3 (.I(_2562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8470__I (.I(_2566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7799__A1 (.I(_2566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7726__A1 (.I(_2566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7307__B (.I(_2566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7383__A1 (.I(_2569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7357__A1 (.I(_2569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7310__A2 (.I(_2569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7691__I (.I(_2574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7450__A2 (.I(_2574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7366__C (.I(_2574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7315__B (.I(_2574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7316__C (.I(_2575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7318__C (.I(_2577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7624__A2 (.I(_2581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7529__A2 (.I(_2581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7477__A2 (.I(_2581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7371__A1 (.I(_2581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8126__A2 (.I(_2582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8086__A1 (.I(_2582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8048__A1 (.I(_2582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7368__A1 (.I(_2582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7622__A2 (.I(_2583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7527__A2 (.I(_2583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7416__A2 (.I(_2583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7368__A2 (.I(_2583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8313__A1 (.I(_2584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8295__A1 (.I(_2584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7673__A1 (.I(_2584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7326__I (.I(_2584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8283__A1 (.I(_2585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8175__A2 (.I(_2585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7458__I (.I(_2585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7327__I (.I(_2585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8320__A2 (.I(_2586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8207__A1 (.I(_2586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8095__A1 (.I(_2586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7328__I (.I(_2586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7704__A1 (.I(_2587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7617__A1 (.I(_2587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7462__A2 (.I(_2587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7332__A1 (.I(_2587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8057__A2 (.I(_2590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7332__A2 (.I(_2590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7369__A1 (.I(_2592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7344__A1 (.I(_2592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7340__A1 (.I(_2592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7334__A1 (.I(_2592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8345__B2 (.I(_2595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8290__B2 (.I(_2595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7337__I (.I(_2595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8433__A1 (.I(_2597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8365__B2 (.I(_2597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7781__A2 (.I(_2597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7339__A2 (.I(_2597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7346__A2 (.I(_2598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7362__B1 (.I(_2599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7345__A2 (.I(_2599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7895__B (.I(_2600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7641__A1 (.I(_2600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7515__A1 (.I(_2600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7344__B (.I(_2600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7611__A1 (.I(_2601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7568__A2 (.I(_2601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7468__A2 (.I(_2601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7343__A1 (.I(_2601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8620__A2 (.I(_2606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8565__C2 (.I(_2606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7664__A1 (.I(_2606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7367__B2 (.I(_2606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7690__A1 (.I(_2607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7606__B2 (.I(_2607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7558__C (.I(_2607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7366__A1 (.I(_2607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7677__I (.I(_2612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7656__B (.I(_2612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7397__C (.I(_2612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7354__C (.I(_2612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7362__A2 (.I(_2619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7804__B2 (.I(_2620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7597__A1 (.I(_2620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7441__I (.I(_2620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7362__B2 (.I(_2620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7367__C (.I(_2625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7914__C (.I(_2629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7905__C (.I(_2629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7873__C (.I(_2629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7371__C (.I(_2629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7418__A1 (.I(_2630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7410__A1 (.I(_2630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7403__A1 (.I(_2630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7374__A1 (.I(_2630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7411__A2 (.I(_2632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7400__A2 (.I(_2632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8786__A2 (.I(_2639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7409__A2 (.I(_2639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7397__A1 (.I(_2639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7389__A1 (.I(_2639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7400__C (.I(_2657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7414__A2 (.I(_2658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8095__A2 (.I(_2660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7404__A2 (.I(_2660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8129__A1 (.I(_2663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8096__A1 (.I(_2663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8094__A1 (.I(_2663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7406__I (.I(_2663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8124__A1 (.I(_2664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8105__A1 (.I(_2664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8087__A1 (.I(_2664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7407__A1 (.I(_2664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7413__A1 (.I(_2665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8093__A2 (.I(_2666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7695__A1 (.I(_2666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7612__A1 (.I(_2666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7411__A1 (.I(_2666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7416__B1 (.I(_2672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7871__A1 (.I(_2673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7745__I (.I(_2673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7621__B (.I(_2673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7416__B2 (.I(_2673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7623__B (.I(_2675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7527__C (.I(_2675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7476__B (.I(_2675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7418__A2 (.I(_2675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7804__A1 (.I(_2678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7730__A1 (.I(_2678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7658__B (.I(_2678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7442__A1 (.I(_2678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7491__A2 (.I(_2679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7490__A2 (.I(_2679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7423__A2 (.I(_2679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7827__A1 (.I(_2686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7758__B2 (.I(_2686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7678__A1 (.I(_2686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7430__B (.I(_2686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7435__A2 (.I(_2691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8550__I (.I(_2693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8517__I (.I(_2693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7585__C (.I(_2693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7437__C (.I(_2693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7442__A2 (.I(_2695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7469__A2 (.I(_2697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7442__B1 (.I(_2697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7762__A1 (.I(_2698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7682__A1 (.I(_2698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7487__A2 (.I(_2698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7442__B2 (.I(_2698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7831__C (.I(_2700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7763__C (.I(_2700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7683__C (.I(_2700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7451__A1 (.I(_2700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7518__C (.I(_2704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7459__B (.I(_2704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7448__B (.I(_2704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7451__A2 (.I(_2706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7528__A1 (.I(_2707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7451__B (.I(_2707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7476__A1 (.I(_2709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8139__A1 (.I(_2710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8130__A1 (.I(_2710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7481__A1 (.I(_2710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7475__A1 (.I(_2710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7485__A1 (.I(_2711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7462__A1 (.I(_2711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8330__I (.I(_2712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8298__A1 (.I(_2712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7865__A2 (.I(_2712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7457__A1 (.I(_2712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8385__A1 (.I(_2713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8099__A1 (.I(_2713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7457__A2 (.I(_2713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7705__B (.I(_2714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7618__B2 (.I(_2714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7522__B (.I(_2714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7462__B (.I(_2714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7996__A1 (.I(_2715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7616__A2 (.I(_2715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7565__S (.I(_2715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7461__A1 (.I(_2715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8141__A2 (.I(_2717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7461__A2 (.I(_2717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7844__B (.I(_2721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7811__B (.I(_2721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7737__B (.I(_2721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7465__I (.I(_2721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8410__A2 (.I(_2722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7569__A1 (.I(_2722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7516__A1 (.I(_2722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7469__A1 (.I(_2722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8297__A2 (.I(_2723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8223__A1 (.I(_2723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7568__B (.I(_2723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7468__B (.I(_2723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8351__A1 (.I(_2728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7784__A2 (.I(_2728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7707__I (.I(_2728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7472__I (.I(_2728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7644__A2 (.I(_2729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7571__B2 (.I(_2729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7524__B2 (.I(_2729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7473__B2 (.I(_2729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8191__B (.I(_2731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8160__B (.I(_2731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8085__I (.I(_2731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7475__B2 (.I(_2731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7700__A1 (.I(_2735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7613__A1 (.I(_2735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7563__A1 (.I(_2735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7483__A1 (.I(_2735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7498__A1 (.I(_2736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7491__A1 (.I(_2736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7490__A1 (.I(_2736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7481__A2 (.I(_2736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7537__A2 (.I(_2738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7483__A2 (.I(_2738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7509__A2 (.I(_2739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7529__A1 (.I(_2740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7522__A1 (.I(_2740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7513__A1 (.I(_2740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7486__A1 (.I(_2740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7516__A2 (.I(_2742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7487__A3 (.I(_2742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7799__B2 (.I(_2744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7726__B2 (.I(_2744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7547__B (.I(_2744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7497__A1 (.I(_2744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7674__A1 (.I(_2759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7504__I (.I(_2759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8598__A1 (.I(_2762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8570__A1 (.I(_2762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8471__A1 (.I(_2762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7507__B (.I(_2762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7509__C (.I(_2764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7602__A1 (.I(_2766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7536__A1 (.I(_2766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7517__A1 (.I(_2766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7511__I (.I(_2766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8215__A1 (.I(_2767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8175__A1 (.I(_2767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8165__A1 (.I(_2767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7524__A1 (.I(_2767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7984__A1 (.I(_2768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7843__A1 (.I(_2768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7779__A2 (.I(_2768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7513__A2 (.I(_2768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7537__A1 (.I(_2773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7520__A1 (.I(_2773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7700__A2 (.I(_2775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7613__A2 (.I(_2775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7563__A2 (.I(_2775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7520__A2 (.I(_2775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8423__C (.I(_2781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8194__I (.I(_2781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7988__I (.I(_2781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7526__I (.I(_2781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8464__A1 (.I(_2782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8302__A1 (.I(_2782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8230__A1 (.I(_2782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7527__B2 (.I(_2782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7528__B (.I(_2783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8233__A1 (.I(_2789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8215__B (.I(_2789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8196__A1 (.I(_2789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7573__A1 (.I(_2789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7700__A3 (.I(_2790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7601__A2 (.I(_2790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7539__A1 (.I(_2790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7560__A2 (.I(_2794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7831__A1 (.I(_2795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7763__A1 (.I(_2795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7683__A1 (.I(_2795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7558__A1 (.I(_2795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7558__A2 (.I(_2807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7830__A1 (.I(_2808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7730__B2 (.I(_2808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7659__A1 (.I(_2808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7557__A1 (.I(_2808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7576__A1 (.I(_2809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7568__A1 (.I(_2809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7565__I0 (.I(_2809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7556__A1 (.I(_2809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7569__A2 (.I(_2811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7557__A2 (.I(_2811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7560__B (.I(_2813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8600__C (.I(_2814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7816__A1 (.I(_2814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7744__A1 (.I(_2814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7560__C (.I(_2814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8447__B (.I(_2816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8354__A1 (.I(_2816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8121__C (.I(_2816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7572__A1 (.I(_2816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7614__A2 (.I(_2817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7564__A1 (.I(_2817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8498__A1 (.I(_2821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7844__A2 (.I(_2821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7640__A2 (.I(_2821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7567__A1 (.I(_2821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7568__C (.I(_2822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7570__B (.I(_2824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7624__A1 (.I(_2832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7616__A1 (.I(_2832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7608__A1 (.I(_2832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7596__A1 (.I(_2832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7766__B (.I(_2840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7715__A2 (.I(_2840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7645__I (.I(_2840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7587__A1 (.I(_2840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7593__A2 (.I(_2845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7606__A1 (.I(_2848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7612__A2 (.I(_2850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7597__A2 (.I(_2850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7606__B1 (.I(_2859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7621__A1 (.I(_2860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8300__A1 (.I(_2861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8228__C (.I(_2861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7848__B2 (.I(_2861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7620__A2 (.I(_2861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8137__A2 (.I(_2863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7984__A3 (.I(_2863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7777__I (.I(_2863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7610__I (.I(_2863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8173__A1 (.I(_2864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8138__A1 (.I(_2864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7694__B (.I(_2864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7611__B (.I(_2864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8250__A2 (.I(_2869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7617__A2 (.I(_2869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7618__B1 (.I(_2871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7620__A3 (.I(_2872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8309__A1 (.I(_2879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7665__A1 (.I(_2879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7644__A1 (.I(_2879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7642__A1 (.I(_2879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7699__A1 (.I(_2882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7687__C (.I(_2882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7660__B (.I(_2882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7630__B (.I(_2882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8283__A2 (.I(_2884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7635__A2 (.I(_2884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7847__A1 (.I(_2886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7814__A1 (.I(_2886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7741__A1 (.I(_2886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7634__B (.I(_2886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7659__A2 (.I(_2890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7641__A2 (.I(_2890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8318__A2 (.I(_2891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8316__A1 (.I(_2891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8003__A2 (.I(_2891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7640__B (.I(_2891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8294__A1 (.I(_2898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7716__A2 (.I(_2898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7653__A1 (.I(_2898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7646__A1 (.I(_2898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8383__A1 (.I(_2903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7734__A1 (.I(_2903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7656__A1 (.I(_2903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7651__A1 (.I(_2903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7753__A1 (.I(_2907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7722__A1 (.I(_2907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7675__A1 (.I(_2907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7655__A3 (.I(_2907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7663__A1 (.I(_2911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7662__A2 (.I(_2914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7664__C (.I(_2916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8551__A1 (.I(_2929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7827__B2 (.I(_2929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7758__A1 (.I(_2929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7678__B2 (.I(_2929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7683__A2 (.I(_2930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7712__A1 (.I(_2931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7705__A1 (.I(_2931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7693__A1 (.I(_2931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7681__A1 (.I(_2931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7695__A2 (.I(_2933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7682__A2 (.I(_2933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7710__A1 (.I(_2935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7702__A1 (.I(_2936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7701__B (.I(_2936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7689__A1 (.I(_2936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7688__A1 (.I(_2936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7768__A1 (.I(_2940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7717__A2 (.I(_2940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7692__A1 (.I(_2940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7690__A2 (.I(_2941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8475__I (.I(_2943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7838__B (.I(_2943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7771__B (.I(_2943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7692__B (.I(_2943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8329__A2 (.I(_2955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8321__A2 (.I(_2955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7704__A2 (.I(_2955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7705__C (.I(_2956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7848__A2 (.I(_2959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7815__A2 (.I(_2959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7743__A2 (.I(_2959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7708__B2 (.I(_2959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8855__A1 (.I(_2961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7816__B2 (.I(_2961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7744__B2 (.I(_2961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7710__B2 (.I(_2961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8341__A1 (.I(_2965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7746__A1 (.I(_2965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7743__A1 (.I(_2965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7740__A1 (.I(_2965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7731__A2 (.I(_2969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8349__A1 (.I(_2970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7736__A2 (.I(_2970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7720__I (.I(_2970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8366__A1 (.I(_2972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8348__A1 (.I(_2972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7724__A1 (.I(_2972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7722__C (.I(_2972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7730__A2 (.I(_2977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7747__A1 (.I(_2978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7737__A1 (.I(_2978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7735__A1 (.I(_2978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7729__A1 (.I(_2978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7739__A2 (.I(_2980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7730__B1 (.I(_2980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7731__B (.I(_2981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8342__A2 (.I(_2984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7734__A2 (.I(_2984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8877__A4 (.I(_2989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7845__C (.I(_2989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7812__C (.I(_2989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7739__C (.I(_2989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7740__B (.I(_2990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8782__A1 (.I(_2993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8490__A1 (.I(_2993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7815__B2 (.I(_2993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7743__B2 (.I(_2993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8412__A2 (.I(_2999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8386__A1 (.I(_2999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7792__A1 (.I(_2999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7750__I (.I(_2999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8371__A1 (.I(_3000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8361__A1 (.I(_3000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7787__A1 (.I(_3000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7781__A1 (.I(_3000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7756__A3 (.I(_3002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7753__C (.I(_3002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7823__A2 (.I(_3006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7798__A2 (.I(_3006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7757__B (.I(_3006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7763__A2 (.I(_3008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7789__A1 (.I(_3009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7779__A1 (.I(_3009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7775__A1 (.I(_3009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7761__A1 (.I(_3009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7780__A2 (.I(_3011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7762__A2 (.I(_3011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7786__A1 (.I(_3013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7771__A2 (.I(_3020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8362__A2 (.I(_3024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7776__A2 (.I(_3024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8364__A2 (.I(_3027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8243__A1 (.I(_3027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8092__A1 (.I(_3027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7780__A1 (.I(_3027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7781__B2 (.I(_3030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8442__C (.I(_3033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8372__C (.I(_3033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8007__C (.I(_3033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7784__B2 (.I(_3033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8567__B (.I(_3038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7851__B (.I(_3038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7818__B (.I(_3038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7789__B (.I(_3038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7832__A2 (.I(_3040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7807__A1 (.I(_3040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7794__A1 (.I(_3040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7834__A1 (.I(_3041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7806__B (.I(_3041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7793__B (.I(_3041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7805__A2 (.I(_3043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7810__A2 (.I(_3044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7796__I (.I(_3044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7804__A2 (.I(_3048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7818__A1 (.I(_3049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7811__A1 (.I(_3049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7809__A1 (.I(_3049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7803__A1 (.I(_3049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7812__A2 (.I(_3052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7804__B1 (.I(_3052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7805__B (.I(_3053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7813__B (.I(_3061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8450__A2 (.I(_3068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8431__A1 (.I(_3068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8415__A1 (.I(_3068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7821__I (.I(_3068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8403__A1 (.I(_3069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7850__A1 (.I(_3069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7848__A1 (.I(_3069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7846__A1 (.I(_3069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8177__B2 (.I(_3070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7843__A2 (.I(_3070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7826__A1 (.I(_3070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7824__A1 (.I(_3070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7831__A2 (.I(_3075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7845__A2 (.I(_3077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7830__A2 (.I(_3077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7849__A1 (.I(_3079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7838__A2 (.I(_3085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7846__B (.I(_3093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7869__A2 (.I(_3100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7985__B (.I(_3101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7890__A1 (.I(_3101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7868__A1 (.I(_3101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7876__A2 (.I(_3102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7859__A2 (.I(_3102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7859__A3 (.I(_3104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7867__A2 (.I(_3107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7889__A1 (.I(_3108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7867__A3 (.I(_3108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7866__A3 (.I(_3110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7972__A1 (.I(_3111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7884__A2 (.I(_3111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7865__A3 (.I(_3111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7866__A4 (.I(_3112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7871__B1 (.I(_3117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7876__A3 (.I(_3121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7982__A1 (.I(_3122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7891__A2 (.I(_3122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7982__A2 (.I(_3125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7891__A3 (.I(_3125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7963__A2 (.I(_3126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7881__A2 (.I(_3126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8178__A1 (.I(_3128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8144__C (.I(_3128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8005__I (.I(_3128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7884__A1 (.I(_3128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7884__B (.I(_3129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7885__A4 (.I(_3130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8217__B (.I(_3132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8100__A1 (.I(_3132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7999__I (.I(_3132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7888__A2 (.I(_3132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8802__A1 (.I(_3133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7888__A4 (.I(_3133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7889__A3 (.I(_3134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7892__A2 (.I(_3137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8410__C (.I(_3139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8323__B2 (.I(_3139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7896__A1 (.I(_3139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7895__A1 (.I(_3139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8097__A2 (.I(_3140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7998__A2 (.I(_3140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7896__A3 (.I(_3140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7905__A2 (.I(_3149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7983__A1 (.I(_3155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7911__C (.I(_3155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7918__A1 (.I(_3156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7916__A2 (.I(_3156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7914__A1 (.I(_3156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7913__A2 (.I(_3156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8232__C (.I(_3161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8193__C (.I(_3161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8163__C (.I(_3161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7918__C (.I(_3161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8457__A3 (.I(_3162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8411__C (.I(_3162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8391__B2 (.I(_3162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7922__A2 (.I(_3162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7922__A4 (.I(_3164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7964__S (.I(_3165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7946__I (.I(_3165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7923__I (.I(_3165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7942__S (.I(_3166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7937__S (.I(_3166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7931__A2 (.I(_3166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7930__A1 (.I(_3166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8846__B (.I(_3167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8832__A2 (.I(_3167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7929__A1 (.I(_3167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8797__A1 (.I(_3168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8501__A1 (.I(_3168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8049__A1 (.I(_3168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7926__I (.I(_3168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8841__A1 (.I(_3169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8493__A1 (.I(_3169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8026__C (.I(_3169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7927__I (.I(_3169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8180__B2 (.I(_3170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7949__I (.I(_3170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7940__A1 (.I(_3170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7928__A1 (.I(_3170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8846__A2 (.I(_3171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8832__B1 (.I(_3171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7929__A2 (.I(_3171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7930__A2 (.I(_3172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8875__A1 (.I(_3174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7960__A2 (.I(_3174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7945__A2 (.I(_3174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7936__A1 (.I(_3174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8420__A1 (.I(_3175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8257__A1 (.I(_3175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8068__A1 (.I(_3175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7934__I (.I(_3175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8830__A1 (.I(_3176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8396__A1 (.I(_3176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7951__A2 (.I(_3176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7935__A2 (.I(_3176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8889__A1 (.I(_3178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7937__I0 (.I(_3178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8810__A2 (.I(_3181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7941__A2 (.I(_3181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8871__A2 (.I(_3182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7942__I0 (.I(_3182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8900__A1 (.I(_3184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8885__A1 (.I(_3184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7945__B (.I(_3184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8901__A1 (.I(_3185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8886__A1 (.I(_3185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7947__I0 (.I(_3185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7961__S (.I(_3186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7955__S (.I(_3186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7953__S (.I(_3186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7947__S (.I(_3186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8374__A1 (.I(_3188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8370__A1 (.I(_3188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8324__B2 (.I(_3188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7950__A1 (.I(_3188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8898__A1 (.I(_3191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8883__A1 (.I(_3191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7953__I0 (.I(_3191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8803__B2 (.I(_3194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8445__A1 (.I(_3194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8285__A1 (.I(_3194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7958__I (.I(_3194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8859__A1 (.I(_3195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8809__C (.I(_3195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8331__A1 (.I(_3195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7959__A1 (.I(_3195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8893__A1 (.I(_3196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7960__B (.I(_3196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8895__A1 (.I(_3197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7961__I0 (.I(_3197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7964__I0 (.I(_3199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7968__A2 (.I(_3201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8874__A1 (.I(_3202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8857__A1 (.I(_3202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8549__A1 (.I(_3202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7968__B (.I(_3202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7977__A1 (.I(_3203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7971__A1 (.I(_3203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7971__B (.I(_3204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7977__B1 (.I(_3206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8878__A2 (.I(_3208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7975__A3 (.I(_3208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7980__C (.I(_3212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7983__A2 (.I(_3213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7983__A3 (.I(_3214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7983__A4 (.I(_3215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8035__A2 (.I(_3218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7986__A2 (.I(_3218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8161__I (.I(_3219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8039__I (.I(_3219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7987__I (.I(_3219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8399__C (.I(_3220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8333__C (.I(_3220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8122__C (.I(_3220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8034__A1 (.I(_3220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8303__A1 (.I(_3221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8192__A1 (.I(_3221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8162__A1 (.I(_3221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8033__A2 (.I(_3221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8028__A1 (.I(_3222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7997__A1 (.I(_3222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7993__I1 (.I(_3222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7992__I0 (.I(_3222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7992__S (.I(_3224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8000__A2 (.I(_3227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8000__B (.I(_3231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8458__B (.I(_3232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8392__B (.I(_3232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8255__B2 (.I(_3232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8000__C (.I(_3232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8350__B2 (.I(_3234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8297__B (.I(_3234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8222__B (.I(_3234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8002__I (.I(_3234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8460__A3 (.I(_3235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8394__B2 (.I(_3235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8245__A1 (.I(_3235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8007__A1 (.I(_3235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8007__A2 (.I(_3237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8418__C1 (.I(_3238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8347__A1 (.I(_3238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8299__B2 (.I(_3238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8006__A1 (.I(_3238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8263__A2 (.I(_3241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8201__A2 (.I(_3241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8019__I (.I(_3241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8009__I (.I(_3241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8279__A2 (.I(_3242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8262__A2 (.I(_3242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8075__A2 (.I(_3242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8016__A2 (.I(_3242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8149__I (.I(_3243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8011__I (.I(_3243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8263__B1 (.I(_3244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8203__B1 (.I(_3244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8021__I (.I(_3244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8012__I (.I(_3244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8262__B1 (.I(_3245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8118__B1 (.I(_3245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8115__B1 (.I(_3245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8016__B1 (.I(_3245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8203__A2 (.I(_3246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8199__A2 (.I(_3246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8070__I (.I(_3246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8014__A2 (.I(_3246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8023__A2 (.I(_3249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8815__A1 (.I(_3250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8265__A2 (.I(_3250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8114__A2 (.I(_3250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8020__A2 (.I(_3250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8279__B1 (.I(_3251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8265__B1 (.I(_3251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8114__B1 (.I(_3251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8020__B1 (.I(_3251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8183__A2 (.I(_3252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8118__A2 (.I(_3252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8115__A2 (.I(_3252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8020__C1 (.I(_3252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8023__B1 (.I(_3253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8155__B1 (.I(_3254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8075__B1 (.I(_3254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8073__B1 (.I(_3254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8022__A2 (.I(_3254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8487__A2 (.I(_3256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8032__B1 (.I(_3256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8811__A1 (.I(_3258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8301__B2 (.I(_3258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8121__B2 (.I(_3258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8032__B2 (.I(_3258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8256__A1 (.I(_3260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8226__A1 (.I(_3260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8145__B (.I(_3260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8028__A2 (.I(_3260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8268__I (.I(_3263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8041__I (.I(_3263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8031__C (.I(_3263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8033__B (.I(_3265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8400__I (.I(_3268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8081__I (.I(_3268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8036__I (.I(_3268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8334__A2 (.I(_3269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8271__A2 (.I(_3269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8124__A2 (.I(_3269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8037__A2 (.I(_3269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8465__C (.I(_3271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8448__C (.I(_3271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8303__B (.I(_3271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8040__I (.I(_3271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8232__A2 (.I(_3272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8193__A2 (.I(_3272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8163__A2 (.I(_3272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8084__A2 (.I(_3272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8425__A1 (.I(_3273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8270__A1 (.I(_3273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8082__A1 (.I(_3273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8080__B (.I(_3273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8062__A2 (.I(_3274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8043__I (.I(_3274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8418__B2 (.I(_3277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8180__A1 (.I(_3277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8146__A1 (.I(_3277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8046__I (.I(_3277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8442__B2 (.I(_3278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8372__B2 (.I(_3278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8106__A1 (.I(_3278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8067__A1 (.I(_3278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8104__A2 (.I(_3279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8048__A2 (.I(_3279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8350__A1 (.I(_3281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8286__I (.I(_3281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8224__A1 (.I(_3281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8050__I (.I(_3281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8255__A1 (.I(_3282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8128__I (.I(_3282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8106__B2 (.I(_3282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8067__B2 (.I(_3282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8056__A2 (.I(_3286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8344__A1 (.I(_3287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8056__A3 (.I(_3287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8065__A1 (.I(_3288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8058__B (.I(_3289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8068__A2 (.I(_3290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8059__A2 (.I(_3290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8064__A2 (.I(_3291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8177__A2 (.I(_3292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8143__A2 (.I(_3292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8098__A2 (.I(_3292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8063__A2 (.I(_3292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8290__A2 (.I(_3293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8140__I (.I(_3293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8063__B1 (.I(_3293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8066__A2 (.I(_3297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8069__B (.I(_3300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8261__A2 (.I(_3302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8154__A2 (.I(_3302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8074__A2 (.I(_3302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8072__A2 (.I(_3302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8815__A2 (.I(_3303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8261__B1 (.I(_3303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8074__B1 (.I(_3303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8072__B1 (.I(_3303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8520__A2 (.I(_3308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8077__A2 (.I(_3308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8821__B (.I(_3310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8527__C (.I(_3310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8258__A1 (.I(_3310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8079__C (.I(_3310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8354__B (.I(_3313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8270__C (.I(_3313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8230__B (.I(_3313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8082__C (.I(_3313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8465__A1 (.I(_3316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8399__A1 (.I(_3316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8333__A1 (.I(_3316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8122__A1 (.I(_3316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8092__A2 (.I(_3322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8093__B (.I(_3323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8101__A2 (.I(_3324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8110__A2 (.I(_3326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8099__A2 (.I(_3326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8121__A2 (.I(_3327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8109__A2 (.I(_3327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8106__B1 (.I(_3327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8098__B1 (.I(_3327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8102__A2 (.I(_3332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8111__A1 (.I(_3334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8463__B2 (.I(_3339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8443__A1 (.I(_3339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8375__A1 (.I(_3339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8110__A1 (.I(_3339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8111__B (.I(_3341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8499__A3 (.I(_3343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8198__I (.I(_3343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8148__I (.I(_3343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8113__I (.I(_3343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8829__A1 (.I(_3344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8423__B1 (.I(_3344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8301__A1 (.I(_3344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8121__A1 (.I(_3344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8184__B1 (.I(_3347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8182__B1 (.I(_3347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8151__B1 (.I(_3347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8117__B1 (.I(_3347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8544__A2 (.I(_3350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8120__I (.I(_3350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8121__B1 (.I(_3351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8466__B (.I(_3354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8401__B (.I(_3354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8334__B (.I(_3354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8124__B (.I(_3354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8162__A2 (.I(_3357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8159__A2 (.I(_3357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8147__A2 (.I(_3357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8214__A4 (.I(_3359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8167__A2 (.I(_3359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8130__A2 (.I(_3359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8146__A2 (.I(_3360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8138__A2 (.I(_3366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8145__A1 (.I(_3368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8158__A2 (.I(_3369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8144__A2 (.I(_3369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8789__B (.I(_3370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8252__B1 (.I(_3370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8177__B1 (.I(_3370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8143__B1 (.I(_3370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8157__A2 (.I(_3372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8143__C1 (.I(_3372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8144__B (.I(_3373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8146__B (.I(_3375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8785__I (.I(_3378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8267__A1 (.I(_3378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8190__A1 (.I(_3378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8159__A1 (.I(_3378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8200__B1 (.I(_3379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8185__B1 (.I(_3379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8183__B1 (.I(_3379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8150__I (.I(_3379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8684__A2 (.I(_3380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8281__B1 (.I(_3380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8278__B1 (.I(_3380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8153__B1 (.I(_3380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8156__A2 (.I(_3383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8559__B1 (.I(_3386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8159__B1 (.I(_3386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8159__C (.I(_3388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8378__B (.I(_3391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8273__I (.I(_3391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8192__C (.I(_3391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8162__C (.I(_3391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8174__A2 (.I(_3394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8166__I (.I(_3394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8192__A2 (.I(_3395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8190__A2 (.I(_3395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8187__A2 (.I(_3395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8181__A2 (.I(_3395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8180__A2 (.I(_3397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8173__A2 (.I(_3400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8179__A1 (.I(_3402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8188__A2 (.I(_3405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8177__C1 (.I(_3405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8180__B1 (.I(_3408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8575__A2 (.I(_3415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8190__B1 (.I(_3415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8189__A2 (.I(_3417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8448__A1 (.I(_3422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8360__A1 (.I(_3422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8355__A1 (.I(_3422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8231__A1 (.I(_3422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8211__A1 (.I(_3424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8197__I (.I(_3424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8231__A2 (.I(_3425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8229__A2 (.I(_3425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8226__A2 (.I(_3425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8224__A2 (.I(_3425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8824__A1 (.I(_3426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8446__B1 (.I(_3426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8353__B1 (.I(_3426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8229__A1 (.I(_3426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8588__B1 (.I(_3432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8229__B1 (.I(_3432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8446__A1 (.I(_3433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8423__A1 (.I(_3433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8353__A1 (.I(_3433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8229__B2 (.I(_3433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8225__A2 (.I(_3435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8212__A3 (.I(_3435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8459__A2 (.I(_3436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8390__A1 (.I(_3436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8211__A2 (.I(_3436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8211__B1 (.I(_3438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8455__A1 (.I(_3441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8346__A1 (.I(_3441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8293__A1 (.I(_3441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8216__A1 (.I(_3441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8217__A2 (.I(_3444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8240__A2 (.I(_3448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8221__A3 (.I(_3448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8223__A2 (.I(_3449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8224__B (.I(_3451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8421__C (.I(_3455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8257__C (.I(_3455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8245__B (.I(_3455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8228__B2 (.I(_3455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8229__C (.I(_3456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8253__A2 (.I(_3461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8235__I (.I(_3461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8270__A2 (.I(_3462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8267__A2 (.I(_3462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8256__A2 (.I(_3462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8255__A2 (.I(_3462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8460__A2 (.I(_3463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8457__A2 (.I(_3463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8436__A2 (.I(_3463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8244__A2 (.I(_3463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8242__A2 (.I(_3467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8241__A2 (.I(_3467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8244__B1 (.I(_3468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8245__A2 (.I(_3471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8453__A2 (.I(_3473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8391__A1 (.I(_3473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8310__A2 (.I(_3473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8254__A1 (.I(_3473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8254__A2 (.I(_3474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8345__A1 (.I(_3475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8321__C (.I(_3475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8292__A1 (.I(_3475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8251__A1 (.I(_3475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8257__A2 (.I(_3477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8251__A2 (.I(_3477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8253__C (.I(_3479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8270__B1 (.I(_3486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8601__A2 (.I(_3493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8269__A2 (.I(_3493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8271__B (.I(_3497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8290__B1 (.I(_3501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8276__I (.I(_3501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8303__A2 (.I(_3502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8301__A2 (.I(_3502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8299__A2 (.I(_3502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8285__A2 (.I(_3502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8617__B1 (.I(_3508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8301__B1 (.I(_3508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8442__A1 (.I(_3512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8418__A1 (.I(_3512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8312__I (.I(_3512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8299__A1 (.I(_3512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8309__A2 (.I(_3513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8308__A3 (.I(_3513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8288__A2 (.I(_3513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8788__A2 (.I(_3515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8291__A2 (.I(_3515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8296__A2 (.I(_3521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8298__A2 (.I(_3523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8301__C (.I(_3526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8322__A2 (.I(_3531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8307__I (.I(_3531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8333__A2 (.I(_3532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8331__A2 (.I(_3532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8327__B2 (.I(_3532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8324__A2 (.I(_3532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8459__A1 (.I(_3537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8394__A1 (.I(_3537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8372__A1 (.I(_3537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8324__A1 (.I(_3537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8366__A4 (.I(_3540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8348__A3 (.I(_3540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8316__A2 (.I(_3540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8322__C (.I(_3546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8324__B1 (.I(_3548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8331__B (.I(_3554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8463__C (.I(_3555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8419__A1 (.I(_3555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8375__B (.I(_3555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8331__C (.I(_3555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8345__B1 (.I(_3561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8338__I (.I(_3561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8355__A2 (.I(_3562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8353__B2 (.I(_3562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8351__B1 (.I(_3562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8350__A2 (.I(_3562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8412__A3 (.I(_3563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8386__A2 (.I(_3563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8371__A2 (.I(_3563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8346__A2 (.I(_3563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8345__C (.I(_3568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8350__B1 (.I(_3573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8353__C (.I(_3576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8365__B1 (.I(_3581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8359__I (.I(_3581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8374__A2 (.I(_3585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8365__A2 (.I(_3585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8365__C (.I(_3587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8437__A3 (.I(_3590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8393__A2 (.I(_3590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8369__B1 (.I(_3590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8369__B2 (.I(_3591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8373__A1 (.I(_3593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8377__A1 (.I(_3597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8450__A4 (.I(_3602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8431__A3 (.I(_3602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8404__A2 (.I(_3602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8381__A2 (.I(_3602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8398__A1 (.I(_3606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8385__A2 (.I(_3606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8391__B1 (.I(_3611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8394__B1 (.I(_3615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8466__A2 (.I(_3622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8429__A2 (.I(_3622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8425__C (.I(_3622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8401__A2 (.I(_3622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8427__A1 (.I(_3624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8425__A2 (.I(_3627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8423__B2 (.I(_3627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8420__A2 (.I(_3627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8418__A2 (.I(_3627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8422__A1 (.I(_3632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8440__A2 (.I(_3633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8413__A2 (.I(_3633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8421__A2 (.I(_3636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8417__A2 (.I(_3636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8424__A1 (.I(_3643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8890__B (.I(_3647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8887__B (.I(_3647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8884__B (.I(_3647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8427__B (.I(_3647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8902__B (.I(_3648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8899__B (.I(_3648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8896__B (.I(_3648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8449__A1 (.I(_3648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8448__A2 (.I(_3652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8446__B2 (.I(_3652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8433__A2 (.I(_3652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8444__A2 (.I(_3654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8435__B1 (.I(_3654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8443__A2 (.I(_3658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8445__A2 (.I(_3659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8442__A2 (.I(_3659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8465__A2 (.I(_3670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8463__B1 (.I(_3670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8462__B2 (.I(_3670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8459__B (.I(_3670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8614__A1 (.I(_3687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8613__C (.I(_3687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8600__A1 (.I(_3687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8476__A1 (.I(_3687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8584__A1 (.I(_3688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8536__A1 (.I(_3688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8516__A1 (.I(_3688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8472__A1 (.I(_3688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8585__C (.I(_3693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8537__C (.I(_3693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8519__C (.I(_3693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8476__C (.I(_3693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8511__A1 (.I(_3694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8847__B1 (.I(_3695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8607__B1 (.I(_3695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8563__B1 (.I(_3695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8478__A2 (.I(_3695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8521__I (.I(_3697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8480__I (.I(_3697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8800__A1 (.I(_3700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8586__A2 (.I(_3700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8557__I (.I(_3700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8483__I (.I(_3700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8604__A2 (.I(_3701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8603__A2 (.I(_3701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8540__A2 (.I(_3701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8484__A2 (.I(_3701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8487__B (.I(_3704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8488__A3 (.I(_3705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8492__C (.I(_3709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8497__A2 (.I(_3714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8508__A3 (.I(_3716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8507__A2 (.I(_3717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8506__A2 (.I(_3723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8507__A4 (.I(_3724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8592__A1 (.I(_3726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8580__B (.I(_3726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8512__I (.I(_3726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8509__I (.I(_3726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8621__A2 (.I(_3727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8569__A2 (.I(_3727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8530__C (.I(_3727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8510__C (.I(_3727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8619__C (.I(_3730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8547__B (.I(_3730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8534__I (.I(_3730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8513__I (.I(_3730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8531__A1 (.I(_3736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8525__A1 (.I(_3737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8527__B1 (.I(_3742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8527__B2 (.I(_3743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8530__B1 (.I(_3744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8548__B1 (.I(_3753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8620__B1 (.I(_3755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8608__B1 (.I(_3755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8564__A1 (.I(_3755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8546__B1 (.I(_3755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8544__B (.I(_3759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8545__C (.I(_3760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8546__B2 (.I(_3761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8554__A2 (.I(_3768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8843__A1 (.I(_3772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8616__A2 (.I(_3772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8574__A2 (.I(_3772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8558__A2 (.I(_3772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8564__A2 (.I(_3776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8847__A2 (.I(_3777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8836__A2 (.I(_3777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8607__A2 (.I(_3777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8563__A2 (.I(_3777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8566__A2 (.I(_3779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8581__B2 (.I(_3786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8579__B1 (.I(_3791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8580__C (.I(_3793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8595__A1 (.I(_3798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8590__A1 (.I(_3800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8860__A1 (.I(_3802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8590__B (.I(_3802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8591__A2 (.I(_3803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8592__A2 (.I(_3804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8609__B (.I(_3812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8606__A1 (.I(_3813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8606__A2 (.I(_3817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8607__C (.I(_3818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8608__B2 (.I(_3819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8614__C (.I(_3824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8622__A1 (.I(_3825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8620__B2 (.I(_3829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8635__I (.I(_3833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8634__I (.I(_3833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8625__I (.I(_3833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8624__I (.I(_3833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8642__A2 (.I(_3841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8640__A2 (.I(_3841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8638__A2 (.I(_3841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8636__A2 (.I(_3841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8650__I (.I(_3846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8645__I (.I(_3846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8661__A2 (.I(_3847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8659__A2 (.I(_3847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8647__I (.I(_3847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8646__I (.I(_3847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8656__A2 (.I(_3848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8654__A2 (.I(_3848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8652__A2 (.I(_3848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8649__A2 (.I(_3848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8662__A2 (.I(_3849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8660__A2 (.I(_3849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8658__A2 (.I(_3849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8648__A2 (.I(_3849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8657__A2 (.I(_3851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8655__A2 (.I(_3851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8653__A2 (.I(_3851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8651__A2 (.I(_3851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8675__I (.I(_3858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8674__I (.I(_3858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8665__I (.I(_3858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8664__I (.I(_3858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8682__A2 (.I(_3866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8680__A2 (.I(_3866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8678__A2 (.I(_3866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8676__A2 (.I(_3866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8701__A2 (.I(_3872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8699__A2 (.I(_3872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8687__I (.I(_3872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8686__I (.I(_3872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8696__A2 (.I(_3873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8694__A2 (.I(_3873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8692__A2 (.I(_3873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8689__A2 (.I(_3873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8702__A2 (.I(_3874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8700__A2 (.I(_3874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8698__A2 (.I(_3874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8688__A2 (.I(_3874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8697__A2 (.I(_3876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8695__A2 (.I(_3876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8693__A2 (.I(_3876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8691__A2 (.I(_3876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8733__A2 (.I(_3883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8731__A2 (.I(_3883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8721__A2 (.I(_3883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8710__A2 (.I(_3883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8736__A2 (.I(_3884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8713__I (.I(_3884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8707__A2 (.I(_3884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8705__I (.I(_3884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8728__B1 (.I(_3890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8722__A2 (.I(_3890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8717__A2 (.I(_3890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8712__A2 (.I(_3890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8728__A2 (.I(_3893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8723__B1 (.I(_3893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8718__B1 (.I(_3893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8715__B1 (.I(_3893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8753__A1 (.I(_3901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8746__A1 (.I(_3901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8743__A1 (.I(_3901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8727__A1 (.I(_3901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8759__A2 (.I(_3906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8756__A2 (.I(_3906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8749__A2 (.I(_3906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8739__A2 (.I(_3906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8755__B1 (.I(_3909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8750__B1 (.I(_3909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8748__B1 (.I(_3909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8738__B1 (.I(_3909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8752__A2 (.I(_3911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8750__A2 (.I(_3911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8745__A2 (.I(_3911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8742__A2 (.I(_3911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8757__A2 (.I(_3912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8752__B1 (.I(_3912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8745__B1 (.I(_3912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8742__B1 (.I(_3912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8772__I (.I(_3924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8771__I (.I(_3924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8762__I (.I(_3924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8761__I (.I(_3924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8833__B2 (.I(_3939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8831__A2 (.I(_3939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8810__C (.I(_3939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8804__A1 (.I(_3939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8866__B1 (.I(_3940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8804__A2 (.I(_3940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8788__B1 (.I(_3941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8803__B1 (.I(_3942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8792__A1 (.I(_3943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8792__A2 (.I(_3944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8792__B (.I(_3945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8841__A2 (.I(_3952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8799__A1 (.I(_3952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8829__B (.I(_3957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8824__B (.I(_3957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8804__B (.I(_3957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8817__A2 (.I(_3959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8816__A1 (.I(_3959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8808__A1 (.I(_3959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8807__A2 (.I(_3959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8822__A2 (.I(_3968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8821__A2 (.I(_3968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8818__A2 (.I(_3968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8816__A2 (.I(_3968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8825__I1 (.I(_3975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8888__A1 (.I(_3976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8824__A2 (.I(_3976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8845__A2 (.I(_3980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8829__A2 (.I(_3980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8833__B1 (.I(_3984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8858__A2 (.I(_3987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8845__A1 (.I(_3987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8839__A4 (.I(_3989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8868__A3 (.I(_3990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8840__I (.I(_3990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8856__A2 (.I(_3996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8849__A1 (.I(_3996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8848__A1 (.I(_3997_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8852__A1 (.I(_4002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8862__A2 (.I(_4011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8865__A2 (.I(_4013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8873__A2 (.I(_4017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8872__B (.I(_4017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8872__A2 (.I(_4018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8891__C (.I(_4025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8878__A3 (.I(_4025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8880__A4 (.I(_4027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8888__A2 (.I(_4028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8885__A2 (.I(_4028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8882__B (.I(_4028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8881__A2 (.I(_4028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8892__A4 (.I(_4036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8900__A2 (.I(_4037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8897__A2 (.I(_4037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8894__B (.I(_4037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8893__A2 (.I(_4037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8901__A2 (.I(_4039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8898__A2 (.I(_4039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8895__A2 (.I(_4039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5876__A1 (.I(_4045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5269__A1 (.I(_4045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5117__A1 (.I(_4045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4452__I (.I(_4045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7045__A1 (.I(_4046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5850__A1 (.I(_4046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5147__A1 (.I(_4046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4453__I (.I(_4046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7925__I (.I(_4047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6106__A1 (.I(_4047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4939__A1 (.I(_4047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4454__I (.I(_4047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8292__B2 (.I(_4048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7880__A1 (.I(_4048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7314__A1 (.I(_4048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4455__I (.I(_4048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8384__C (.I(_4049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8187__A1 (.I(_4049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6292__A1 (.I(_4049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4456__I (.I(_4049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8102__A1 (.I(_4050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8000__A1 (.I(_4050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6404__C (.I(_4050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4457__I (.I(_4050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8894__A1 (.I(_4051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7230__A1 (.I(_4051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7219__A2 (.I(_4051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4664__A1 (.I(_4051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4722__A1 (.I(_4052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4645__I (.I(_4052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4564__A1 (.I(_4052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4459__I (.I(_4052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4711__A2 (.I(_4053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4703__I (.I(_4053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4640__A1 (.I(_4053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4462__A1 (.I(_4053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4639__A1 (.I(_4054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4633__I (.I(_4054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4564__A2 (.I(_4054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4461__I (.I(_4054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5074__I (.I(_4055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4946__A2 (.I(_4055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4656__A1 (.I(_4055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4462__A2 (.I(_4055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8496__A1 (.I(_4057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7994__S (.I(_4057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5148__A1 (.I(_4057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4627__A1 (.I(_4057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4546__S0 (.I(_4058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4537__S0 (.I(_4058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4528__S0 (.I(_4058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4465__I (.I(_4058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4519__S0 (.I(_4059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4499__I (.I(_4059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4493__C (.I(_4059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4466__I (.I(_4059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6110__I (.I(_4060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5057__A1 (.I(_4060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4630__A2 (.I(_4060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4471__S0 (.I(_4060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4568__S1 (.I(_4062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4567__S (.I(_4062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4551__S1 (.I(_4062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4469__I (.I(_4062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4519__S1 (.I(_4063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4502__S (.I(_4063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4488__I (.I(_4063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4470__I (.I(_4063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5114__I (.I(_4064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5107__A1 (.I(_4064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4479__S (.I(_4064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4471__S1 (.I(_4064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4475__A1 (.I(_4065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4551__S0 (.I(_4066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4483__A1 (.I(_4066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4476__A1 (.I(_4066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4473__A1 (.I(_4066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4638__I (.I(_4072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4518__A1 (.I(_4072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4503__A1 (.I(_4072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4480__A1 (.I(_4072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8314__A2 (.I(_4073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8313__A2 (.I(_4073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8295__A2 (.I(_4073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4480__A2 (.I(_4073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6846__A1 (.I(_4075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6704__A1 (.I(_4075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6703__A1 (.I(_4075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4482__I (.I(_4075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6870__A1 (.I(_4076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6758__A1 (.I(_4076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5783__I (.I(_4076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4486__A1 (.I(_4076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4535__A2 (.I(_4078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4525__A2 (.I(_4078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4513__A2 (.I(_4078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4485__I (.I(_4078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5072__I (.I(_4079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4799__I (.I(_4079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4507__A2 (.I(_4079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4486__A2 (.I(_4079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6930__A1 (.I(_4081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6280__I (.I(_4081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5823__A1 (.I(_4081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4590__A1 (.I(_4081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6490__A1 (.I(_4082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5139__I (.I(_4082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4493__A1 (.I(_4082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4489__A1 (.I(_4082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5052__I (.I(_4085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4629__A2 (.I(_4085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4500__A2 (.I(_4085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4492__I (.I(_4085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5056__I (.I(_4086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4779__A2 (.I(_4086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4493__B (.I(_4086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6557__S (.I(_4088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6554__S (.I(_4088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6543__S (.I(_4088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4495__S (.I(_4088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6813__A2 (.I(_4089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6764__A2 (.I(_4089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6668__A2 (.I(_4089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4496__I (.I(_4089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6815__B1 (.I(_4090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6707__A2 (.I(_4090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6633__A2 (.I(_4090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4497__I (.I(_4090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6869__A2 (.I(_4091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6708__B1 (.I(_4091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6669__B1 (.I(_4091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4498__I (.I(_4091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8605__A1 (.I(_4092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6944__A3 (.I(_4092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6916__A2 (.I(_4092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4501__B1 (.I(_4092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5727__I (.I(_4094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5081__A2 (.I(_4094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4501__B2 (.I(_4094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4591__A1 (.I(_4095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4508__A1 (.I(_4095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8294__A2 (.I(_4096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8237__A2 (.I(_4096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4503__A2 (.I(_4096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6869__A1 (.I(_4099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6844__A1 (.I(_4099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6694__A1 (.I(_4099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4506__I (.I(_4099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6808__A1 (.I(_4100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5753__A1 (.I(_4100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5716__I (.I(_4100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4507__A1 (.I(_4100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5731__A2 (.I(_4102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4509__I (.I(_4102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5822__A2 (.I(_4103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5754__A1 (.I(_4103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4587__I (.I(_4103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4510__I (.I(_4103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6689__A1 (.I(_4106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5682__I (.I(_4106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5655__A1 (.I(_4106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4513__A1 (.I(_4106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6656__A1 (.I(_4108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6572__S (.I(_4108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4557__S (.I(_4108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4515__I (.I(_4108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4546__S1 (.I(_4109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4541__S (.I(_4109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4526__S (.I(_4109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4516__I (.I(_4109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4537__S1 (.I(_4110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4536__S (.I(_4110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4528__S1 (.I(_4110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4517__S (.I(_4110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8239__A2 (.I(_4111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8238__A2 (.I(_4111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8221__A2 (.I(_4111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4518__A2 (.I(_4111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4520__A2 (.I(_4113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5677__A1 (.I(_4115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5656__A1 (.I(_4115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4522__I (.I(_4115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5675__B (.I(_4116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5658__A1 (.I(_4116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5650__I (.I(_4116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4574__A1 (.I(_4116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6628__A1 (.I(_4118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6563__A1 (.I(_4118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5582__I (.I(_4118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4525__A1 (.I(_4118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8219__A2 (.I(_4120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8218__A2 (.I(_4120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8171__A2 (.I(_4120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4527__A2 (.I(_4120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4580__A2 (.I(_4121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4530__A2 (.I(_4121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4529__A2 (.I(_4122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4580__A3 (.I(_4123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4530__A3 (.I(_4123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5607__A1 (.I(_4124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4531__I (.I(_4124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5677__A2 (.I(_4125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5608__A1 (.I(_4125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5584__A1 (.I(_4125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4532__I (.I(_4125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6710__A1 (.I(_4127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6635__A1 (.I(_4127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6564__A1 (.I(_4127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4534__I (.I(_4127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6653__A1 (.I(_4128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6582__A1 (.I(_4128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5511__I (.I(_4128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4535__A1 (.I(_4128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4611__A1 (.I(_4129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4605__A1 (.I(_4129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4584__A1 (.I(_4129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4539__A1 (.I(_4129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8132__A2 (.I(_4130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8131__A2 (.I(_4130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4538__A2 (.I(_4130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4538__B1 (.I(_4131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4611__A2 (.I(_4132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4605__A2 (.I(_4132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4584__A2 (.I(_4132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4539__A2 (.I(_4132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6789__A1 (.I(_4134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5540__B2 (.I(_4134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4603__A1 (.I(_4134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4573__A1 (.I(_4134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8134__A2 (.I(_4135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8088__A2 (.I(_4135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4542__A2 (.I(_4135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5535__A1 (.I(_4136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4596__A1 (.I(_4136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4584__A3 (.I(_4136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4543__I (.I(_4136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5435__A1 (.I(_4137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5433__A1 (.I(_4137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4605__A3 (.I(_4137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4549__A1 (.I(_4137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6756__A1 (.I(_4138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6708__A1 (.I(_4138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6559__A1 (.I(_4138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4545__I (.I(_4138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6597__A1 (.I(_4139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6583__B2 (.I(_4139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5436__I (.I(_4139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4547__A1 (.I(_4139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4547__B1 (.I(_4140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5535__A2 (.I(_4141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4596__A2 (.I(_4141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4584__A4 (.I(_4141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4548__I (.I(_4141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5435__A2 (.I(_4142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5433__A2 (.I(_4142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4605__A4 (.I(_4142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4549__A2 (.I(_4142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5486__A1 (.I(_4143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5465__A1 (.I(_4143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4550__I (.I(_4143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5487__A1 (.I(_4144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5382__I (.I(_4144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4620__A1 (.I(_4144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4573__A2 (.I(_4144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4552__A2 (.I(_4145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4614__A1 (.I(_4146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4553__I (.I(_4146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5535__B1 (.I(_4147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5342__A1 (.I(_4147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4583__A1 (.I(_4147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4554__I (.I(_4147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5461__A1 (.I(_4148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5459__A1 (.I(_4148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5354__A1 (.I(_4148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4561__A1 (.I(_4148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6698__A1 (.I(_4150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6566__A1 (.I(_4150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5343__I (.I(_4150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4558__A1 (.I(_4150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8089__A2 (.I(_4151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8052__A2 (.I(_4151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4558__B1 (.I(_4151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4614__A2 (.I(_4152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4559__I (.I(_4152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5535__B2 (.I(_4153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5342__A2 (.I(_4153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4583__A2 (.I(_4153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4560__I (.I(_4153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5461__A2 (.I(_4154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5459__A2 (.I(_4154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5354__A2 (.I(_4154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4561__A2 (.I(_4154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6330__A2 (.I(_4156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5479__A1 (.I(_4156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4619__A1 (.I(_4156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4573__A3 (.I(_4156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4732__A3 (.I(_4157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4722__A2 (.I(_4157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4616__A1 (.I(_4157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4572__A1 (.I(_4157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6522__A1 (.I(_4158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4622__A1 (.I(_4158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4616__A2 (.I(_4158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4572__A2 (.I(_4158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6669__B2 (.I(_4159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6657__A1 (.I(_4159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6545__A2 (.I(_4159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4566__I (.I(_4159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6667__A1 (.I(_4160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6549__A1 (.I(_4160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5178__I (.I(_4160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4569__A1 (.I(_4160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8051__A2 (.I(_4161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8003__A1 (.I(_4161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4569__B1 (.I(_4161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4569__C1 (.I(_4162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5389__I (.I(_4163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4582__I (.I(_4163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4570__I (.I(_4163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5459__B (.I(_4164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5182__A1 (.I(_4164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5176__I1 (.I(_4164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4571__I (.I(_4164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8502__A1 (.I(_4170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5155__A1 (.I(_4170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4577__A2 (.I(_4170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4607__A1 (.I(_4171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4600__A1 (.I(_4171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4592__A1 (.I(_4171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4588__A1 (.I(_4171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5674__A1 (.I(_4172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4579__I (.I(_4172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5606__A1 (.I(_4174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4581__I (.I(_4174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5674__A2 (.I(_4175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5578__A1 (.I(_4175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5544__I (.I(_4175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4585__A2 (.I(_4175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5461__A3 (.I(_4176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5396__A1 (.I(_4176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4599__I (.I(_4176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4583__A3 (.I(_4176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6327__A1 (.I(_4180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4607__A2 (.I(_4180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4592__A2 (.I(_4180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4588__A2 (.I(_4180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5820__A1 (.I(_4181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5755__A1 (.I(_4181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5749__A1 (.I(_4181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4588__A3 (.I(_4181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5814__I (.I(_4184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4627__A2 (.I(_4184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6329__I (.I(_4185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5730__A1 (.I(_4185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4594__A1 (.I(_4185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6364__C1 (.I(_4189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5694__I (.I(_4189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4609__A1 (.I(_4189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4604__A1 (.I(_4189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5462__A1 (.I(_4190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4597__I (.I(_4190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5539__A1 (.I(_4191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5460__A1 (.I(_4191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5430__A1 (.I(_4191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4598__I (.I(_4191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6365__A2 (.I(_4192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5543__I (.I(_4192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4617__A1 (.I(_4192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4602__A1 (.I(_4192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5240__A1 (.I(_4193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5195__A1 (.I(_4193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5190__A1 (.I(_4193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4600__A2 (.I(_4193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8580__A1 (.I(_4198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6888__A1 (.I(_4198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5619__A1 (.I(_4198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4626__A1 (.I(_4198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6328__A3 (.I(_4199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5677__A4 (.I(_4199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4606__A3 (.I(_4199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6931__A1 (.I(_4202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6889__A1 (.I(_4202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5622__I (.I(_4202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4610__I1 (.I(_4202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8594__A1 (.I(_4204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6902__A1 (.I(_4204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5691__A1 (.I(_4204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4626__A2 (.I(_4204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5539__B (.I(_4206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5513__A1 (.I(_4206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5508__A1 (.I(_4206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4613__I (.I(_4206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6368__A2 (.I(_4207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5554__A1 (.I(_4207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5472__I (.I(_4207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4618__A1 (.I(_4207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5397__A1 (.I(_4208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5392__A1 (.I(_4208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5341__A1 (.I(_4208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4615__I (.I(_4208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6368__B1 (.I(_4209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5264__I (.I(_4209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4624__A1 (.I(_4209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4617__A2 (.I(_4209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8565__C1 (.I(_4212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6832__A1 (.I(_4212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5548__A1 (.I(_4212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4625__A1 (.I(_4212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8547__A1 (.I(_4214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6788__A1 (.I(_4214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5476__A1 (.I(_4214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4625__A2 (.I(_4214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6522__A2 (.I(_4215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6365__C1 (.I(_4215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5373__I (.I(_4215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4622__A2 (.I(_4215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5274__A1 (.I(_4216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4625__A3 (.I(_4216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8528__A2 (.I(_4218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6735__A1 (.I(_4218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5380__A1 (.I(_4218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4625__A4 (.I(_4218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8044__A1 (.I(_4221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4628__I (.I(_4221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8049__A2 (.I(_4222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7853__A1 (.I(_4222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5051__A2 (.I(_4222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4664__A2 (.I(_4222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4642__A1 (.I(_4225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4641__A2 (.I(_4225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4870__A1 (.I(_4226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4747__I (.I(_4226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4660__A2 (.I(_4226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4637__A1 (.I(_4226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4945__I (.I(_4228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4655__I (.I(_4228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4639__A2 (.I(_4228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4635__A2 (.I(_4228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5210__A2 (.I(_4230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5172__A1 (.I(_4230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5077__B (.I(_4230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4637__A2 (.I(_4230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4642__A2 (.I(_4231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4694__A1 (.I(_4232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4684__A1 (.I(_4232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4654__I (.I(_4232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4641__A1 (.I(_4232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5054__A2 (.I(_4234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4731__A2 (.I(_4234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4641__A3 (.I(_4234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8793__A1 (.I(_4235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6129__A2 (.I(_4235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4642__B (.I(_4235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7993__S (.I(_4236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5084__A1 (.I(_4236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4643__I (.I(_4236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8049__A3 (.I(_4237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8044__A2 (.I(_4237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7241__A1 (.I(_4237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4664__A3 (.I(_4237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5842__A1 (.I(_4238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4728__A1 (.I(_4238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4699__I (.I(_4238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4646__A1 (.I(_4238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4792__I (.I(_4239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4732__A2 (.I(_4239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4721__A2 (.I(_4239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4646__A2 (.I(_4239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4848__A3 (.I(_4240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4693__A2 (.I(_4240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4685__A2 (.I(_4240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4647__I (.I(_4240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7984__A2 (.I(_4241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7877__A2 (.I(_4241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6161__A1 (.I(_4241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4648__I (.I(_4241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7299__B (.I(_4242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5046__I (.I(_4242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5018__I (.I(_4242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4653__A1 (.I(_4242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6128__A1 (.I(_4243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5854__A1 (.I(_4243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4908__I (.I(_4243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4651__A1 (.I(_4243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6485__A2 (.I(_4245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5858__A2 (.I(_4245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5115__A4 (.I(_4245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4652__I (.I(_4245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6420__A2 (.I(_4246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5865__A1 (.I(_4246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4920__A2 (.I(_4246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4653__A2 (.I(_4246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8798__A1 (.I(_4248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6391__I (.I(_4248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5066__A2 (.I(_4248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4661__A1 (.I(_4248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4825__I (.I(_4249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4724__A1 (.I(_4249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4656__A2 (.I(_4249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4694__A2 (.I(_4250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4684__A2 (.I(_4250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4657__I (.I(_4250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8837__A1 (.I(_4251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5448__A1 (.I(_4251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5206__A2 (.I(_4251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4661__A2 (.I(_4251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6730__A1 (.I(_4253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6112__A1 (.I(_4253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4845__I (.I(_4253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4660__A1 (.I(_4253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4880__A2 (.I(_4255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4811__A2 (.I(_4255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4676__A2 (.I(_4255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4662__I (.I(_4255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7860__A3 (.I(_4256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7049__A1 (.I(_4256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6420__A3 (.I(_4256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4663__A2 (.I(_4256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5084__A2 (.I(_4257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4953__B2 (.I(_4257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4664__A4 (.I(_4257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5166__A1 (.I(_4259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5048__I (.I(_4259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4893__I (.I(_4259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4698__A1 (.I(_4259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5117__A2 (.I(_4261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4972__A2 (.I(_4261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4719__I (.I(_4261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4668__I (.I(_4261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8289__A1 (.I(_4262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7894__A1 (.I(_4262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4736__A2 (.I(_4262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4697__A1 (.I(_4262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7052__A1 (.I(_4265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4900__A2 (.I(_4265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4841__A1 (.I(_4265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4672__A1 (.I(_4265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8047__A2 (.I(_4268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4723__A1 (.I(_4268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4683__I (.I(_4268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4675__I (.I(_4268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4732__A1 (.I(_4269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4730__I (.I(_4269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4711__A1 (.I(_4269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4676__A1 (.I(_4269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7045__A2 (.I(_4270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4918__A4 (.I(_4270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4829__I (.I(_4270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4681__A1 (.I(_4270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4854__I (.I(_4274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4681__A3 (.I(_4274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7875__A2 (.I(_4275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7039__A2 (.I(_4275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5024__B2 (.I(_4275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4695__A2 (.I(_4275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7414__B2 (.I(_4276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7347__I (.I(_4276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7260__A1 (.I(_4276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4692__A1 (.I(_4276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5027__A1 (.I(_4277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4701__I (.I(_4277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4693__A1 (.I(_4277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4686__A1 (.I(_4277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5023__A1 (.I(_4280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4934__I (.I(_4280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4692__A2 (.I(_4280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6506__A2 (.I(_4281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5022__I (.I(_4281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4692__A3 (.I(_4281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8468__I (.I(_4282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5153__A1 (.I(_4282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4918__A2 (.I(_4282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4690__A1 (.I(_4282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7253__A1 (.I(_4283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4879__A2 (.I(_4283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4876__A1 (.I(_4283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4690__A2 (.I(_4283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7232__A2 (.I(_4284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6507__A1 (.I(_4284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4691__A2 (.I(_4284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5860__A1 (.I(_4285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5023__A2 (.I(_4285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4692__A4 (.I(_4285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7984__B (.I(_4286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4695__B (.I(_4286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7049__A2 (.I(_4287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4694__A3 (.I(_4287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5842__A2 (.I(_4288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5014__I (.I(_4288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4695__C (.I(_4288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4697__A2 (.I(_4289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7252__C (.I(_4290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5012__I (.I(_4290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4756__A1 (.I(_4290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4697__B (.I(_4290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6493__A1 (.I(_4293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4775__A1 (.I(_4293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4713__A1 (.I(_4293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4700__I (.I(_4293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8112__A1 (.I(_4294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5007__I (.I(_4294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4773__I (.I(_4294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4707__A1 (.I(_4294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6112__A2 (.I(_4295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4972__A1 (.I(_4295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4811__A1 (.I(_4295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4702__I (.I(_4295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5008__I (.I(_4296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4950__A1 (.I(_4296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4848__A1 (.I(_4296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4706__A1 (.I(_4296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6159__A2 (.I(_4297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5154__A1 (.I(_4297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5081__A1 (.I(_4297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4704__I (.I(_4297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7255__A1 (.I(_4298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6139__A1 (.I(_4298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4790__A1 (.I(_4298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4706__A2 (.I(_4298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8491__A1 (.I(_4299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5447__A2 (.I(_4299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5171__A2 (.I(_4299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4706__A3 (.I(_4299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6156__I (.I(_4300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4707__A2 (.I(_4300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8788__C (.I(_4301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8024__I (.I(_4301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4718__A1 (.I(_4301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4938__A2 (.I(_4304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4711__A3 (.I(_4304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6362__I (.I(_4306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6358__A2 (.I(_4306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4733__A1 (.I(_4306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4713__A2 (.I(_4306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6500__A2 (.I(_4307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5257__A2 (.I(_4307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4714__I (.I(_4307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8800__C (.I(_4308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8492__A2 (.I(_4308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7248__A1 (.I(_4308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4718__A2 (.I(_4308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6495__A2 (.I(_4310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5149__A1 (.I(_4310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5141__A2 (.I(_4310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4717__I (.I(_4310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4770__I (.I(_4311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4736__A1 (.I(_4311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4727__A1 (.I(_4311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4718__B (.I(_4311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5084__C (.I(_4312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4737__A2 (.I(_4312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7336__A2 (.I(_4313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5026__A1 (.I(_4313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4880__A3 (.I(_4313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4720__I (.I(_4313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8495__A2 (.I(_4314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4965__A2 (.I(_4314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4835__I (.I(_4314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4727__A2 (.I(_4314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8491__A2 (.I(_4315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4777__I (.I(_4315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4725__A1 (.I(_4315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6163__A2 (.I(_4317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5029__A2 (.I(_4317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4724__A2 (.I(_4317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8499__A2 (.I(_4318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6331__I (.I(_4318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4725__A2 (.I(_4318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6288__A1 (.I(_4320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6162__A1 (.I(_4320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5034__I (.I(_4320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4727__A3 (.I(_4320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7246__A1 (.I(_4322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5268__A1 (.I(_4322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4729__I (.I(_4322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7227__A1 (.I(_4323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7056__A1 (.I(_4323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4852__I (.I(_4323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4736__A3 (.I(_4323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7336__A1 (.I(_4324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5003__I (.I(_4324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4775__A2 (.I(_4324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4731__A1 (.I(_4324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5267__A2 (.I(_4326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4858__A2 (.I(_4326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4813__A2 (.I(_4326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4733__A2 (.I(_4326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7980__B2 (.I(_4327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4734__A2 (.I(_4327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7246__A2 (.I(_4329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6284__A1 (.I(_4329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6107__B (.I(_4329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4736__A4 (.I(_4329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5118__A2 (.I(_4333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4815__I (.I(_4333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4740__A2 (.I(_4333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7856__A1 (.I(_4334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4741__I (.I(_4334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8505__B (.I(_4335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6173__B (.I(_4335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4824__A2 (.I(_4335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4742__I (.I(_4335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7508__B (.I(_4336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7399__A1 (.I(_4336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7313__A1 (.I(_4336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4746__A1 (.I(_4336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7857__A1 (.I(_4337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7052__A2 (.I(_4337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4886__A1 (.I(_4337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4744__A2 (.I(_4337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6174__A2 (.I(_4338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5133__A1 (.I(_4338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4824__A3 (.I(_4338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4745__I (.I(_4338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7429__I (.I(_4339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7359__C (.I(_4339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7311__I (.I(_4339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4746__A2 (.I(_4339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7236__A2 (.I(_4340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4758__A1 (.I(_4340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7050__A2 (.I(_4341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6429__A1 (.I(_4341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4938__A1 (.I(_4341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4748__I (.I(_4341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6155__I (.I(_4342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4947__A1 (.I(_4342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4891__I (.I(_4342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4757__A1 (.I(_4342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7126__C (.I(_4343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5866__A1 (.I(_4343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4924__I (.I(_4343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4757__A2 (.I(_4343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6165__A2 (.I(_4344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5269__A2 (.I(_4344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5151__A2 (.I(_4344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4751__I (.I(_4344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8061__A1 (.I(_4345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6160__A1 (.I(_4345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4950__A2 (.I(_4345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4752__I (.I(_4345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7244__A2 (.I(_4346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7060__A2 (.I(_4346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4932__I (.I(_4346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4756__A2 (.I(_4346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7253__A2 (.I(_4348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7232__A1 (.I(_4348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6164__A2 (.I(_4348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4755__I (.I(_4348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7901__B2 (.I(_4349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7896__A2 (.I(_4349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5032__A2 (.I(_4349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4756__A3 (.I(_4349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4985__A1 (.I(_4350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4903__A2 (.I(_4350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4757__A3 (.I(_4350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5000__A1 (.I(_4351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4887__A1 (.I(_4351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4827__C (.I(_4351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4758__A2 (.I(_4351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4862__A1 (.I(_4352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4761__A2 (.I(_4352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7228__A1 (.I(_4353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7226__A1 (.I(_4353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7211__A2 (.I(_4353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4760__I (.I(_4353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7213__A1 (.I(_4354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4957__A1 (.I(_4354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4920__A1 (.I(_4354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4761__B (.I(_4354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4833__A1 (.I(_4355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6498__A1 (.I(_4356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5151__A1 (.I(_4356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5108__A1 (.I(_4356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4763__I (.I(_4356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6492__A1 (.I(_4357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6159__A1 (.I(_4357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5326__I (.I(_4357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4764__I (.I(_4357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5864__A1 (.I(_4358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5848__A1 (.I(_4358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5403__I (.I(_4358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4765__I (.I(_4358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8496__B (.I(_4359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6299__A1 (.I(_4359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6170__I (.I(_4359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4766__I (.I(_4359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8252__C (.I(_4360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7044__A1 (.I(_4360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5993__A1 (.I(_4360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4767__I (.I(_4360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8818__B (.I(_4361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8188__A1 (.I(_4361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6137__A2 (.I(_4361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4768__I (.I(_4361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8069__A1 (.I(_4362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7944__A1 (.I(_4362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7620__A1 (.I(_4362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4769__I (.I(_4362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5085__B (.I(_4363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4926__A1 (.I(_4363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4832__A1 (.I(_4363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4814__A1 (.I(_4363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6413__A1 (.I(_4364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5878__A1 (.I(_4364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4853__A1 (.I(_4364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4771__I (.I(_4364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4941__A1 (.I(_4365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4867__I (.I(_4365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4851__A2 (.I(_4365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4772__I (.I(_4365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4992__A2 (.I(_4366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4976__A2 (.I(_4366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4832__A2 (.I(_4366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4814__A2 (.I(_4366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8528__A1 (.I(_4368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8489__C (.I(_4368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8422__B (.I(_4368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4813__A1 (.I(_4368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6324__A2 (.I(_4370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5031__A2 (.I(_4370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4873__A1 (.I(_4370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4810__A1 (.I(_4370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6301__A1 (.I(_4371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6285__C (.I(_4371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5036__A1 (.I(_4371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4809__A1 (.I(_4371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6423__B2 (.I(_4372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6367__A1 (.I(_4372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5060__A1 (.I(_4372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4779__A1 (.I(_4372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5143__A1 (.I(_4373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4780__I (.I(_4373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6492__A2 (.I(_4374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6486__A2 (.I(_4374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6138__I (.I(_4374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4786__A1 (.I(_4374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5181__I (.I(_4375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4782__I (.I(_4375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5656__C (.I(_4376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5340__A2 (.I(_4376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5195__A2 (.I(_4376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4783__I (.I(_4376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5584__C (.I(_4377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5509__A2 (.I(_4377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5430__A2 (.I(_4377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4784__I (.I(_4377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5754__C (.I(_4378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5591__A2 (.I(_4378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5061__I (.I(_4378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4785__I (.I(_4378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5786__C (.I(_4379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5654__A2 (.I(_4379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5059__A2 (.I(_4379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4786__A2 (.I(_4379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5321__A1 (.I(_4380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4938__A3 (.I(_4380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4790__A2 (.I(_4380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5054__A1 (.I(_4381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5027__A2 (.I(_4381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4826__A1 (.I(_4381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4788__A1 (.I(_4381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5081__A4 (.I(_4382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5066__A4 (.I(_4382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5062__A2 (.I(_4382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4789__I (.I(_4382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5520__B (.I(_4383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5457__A1 (.I(_4383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5359__B (.I(_4383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4790__A3 (.I(_4383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7980__A1 (.I(_4384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5067__A1 (.I(_4384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4791__A2 (.I(_4384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8491__A3 (.I(_4385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4809__A2 (.I(_4385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5120__A1 (.I(_4386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5062__A1 (.I(_4386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5058__A1 (.I(_4386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4793__I (.I(_4386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7234__A1 (.I(_4387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6366__A1 (.I(_4387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5066__A1 (.I(_4387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4794__I (.I(_4387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6390__A1 (.I(_4388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4939__A2 (.I(_4388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4806__I (.I(_4388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4805__A1 (.I(_4388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6139__A2 (.I(_4390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5222__A1 (.I(_4390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5214__A1 (.I(_4390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4797__I (.I(_4390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5861__A1 (.I(_4391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5364__A1 (.I(_4391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5070__I (.I(_4391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4805__A2 (.I(_4391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8492__B2 (.I(_4392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7222__A1 (.I(_4392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6251__A2 (.I(_4392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4805__A3 (.I(_4392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6499__A1 (.I(_4393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5270__A1 (.I(_4393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5109__A1 (.I(_4393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4804__A1 (.I(_4393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5354__A3 (.I(_4394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5345__B (.I(_4394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5175__I (.I(_4394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4801__I (.I(_4394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5755__A2 (.I(_4396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5578__A2 (.I(_4396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5053__I (.I(_4396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4803__I (.I(_4396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5787__A2 (.I(_4397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5758__A2 (.I(_4397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4942__I (.I(_4397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4804__A2 (.I(_4397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8891__B (.I(_4398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5328__A1 (.I(_4398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5068__A1 (.I(_4398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4805__A4 (.I(_4398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7966__A2 (.I(_4399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6288__A2 (.I(_4399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4809__B1 (.I(_4399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8499__A1 (.I(_4400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4961__I (.I(_4400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4936__A1 (.I(_4400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4807__I (.I(_4400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7268__A1 (.I(_4401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7046__B (.I(_4401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4874__I (.I(_4401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4808__I (.I(_4401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8866__B2 (.I(_4402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7860__A2 (.I(_4402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6353__I (.I(_4402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4809__B2 (.I(_4402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4810__A2 (.I(_4403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8227__I (.I(_4405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7878__A1 (.I(_4405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7259__A1 (.I(_4405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4812__I (.I(_4405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7847__B2 (.I(_4406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7814__B2 (.I(_4406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7741__B2 (.I(_4406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4813__C (.I(_4406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4814__A3 (.I(_4407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7315__A1 (.I(_4409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4994__I (.I(_4409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4822__A2 (.I(_4409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4816__I (.I(_4409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7838__A1 (.I(_4410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7659__B (.I(_4410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7442__C (.I(_4410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4823__A1 (.I(_4410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7503__A1 (.I(_4411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7294__I (.I(_4411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4837__I (.I(_4411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4819__A2 (.I(_4411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6488__A1 (.I(_4413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5371__A1 (.I(_4413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5127__A1 (.I(_4413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4823__A2 (.I(_4413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6364__A1 (.I(_4414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6354__I (.I(_4414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4986__I (.I(_4414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4821__I (.I(_4414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8284__A2 (.I(_4415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8206__A2 (.I(_4415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7880__A2 (.I(_4415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4822__A1 (.I(_4415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8505__A1 (.I(_4418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4827__A2 (.I(_4418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6169__A2 (.I(_4420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4953__A1 (.I(_4420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4870__A2 (.I(_4420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4827__B (.I(_4420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4828__I (.I(_4421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4833__A3 (.I(_4422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8794__A1 (.I(_4423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8045__A1 (.I(_4423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7893__I (.I(_4423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4830__I (.I(_4423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8788__A1 (.I(_4424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8435__C (.I(_4424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4836__A1 (.I(_4424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4831__I (.I(_4424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8411__A1 (.I(_4425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8369__A1 (.I(_4425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8310__A1 (.I(_4425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4832__A3 (.I(_4425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8363__B (.I(_4428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7895__A2 (.I(_4428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4868__I (.I(_4428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4836__A2 (.I(_4428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8436__B (.I(_4429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8323__A1 (.I(_4429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8101__A1 (.I(_4429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4866__A1 (.I(_4429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7300__A1 (.I(_4430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7290__I (.I(_4430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6173__A1 (.I(_4430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4838__I (.I(_4430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7811__A2 (.I(_4431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7737__A2 (.I(_4431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7467__A1 (.I(_4431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4839__I (.I(_4431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7895__C (.I(_4432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7100__A1 (.I(_4432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4998__B2 (.I(_4432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4851__A1 (.I(_4432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6165__A1 (.I(_4433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4928__I (.I(_4433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4879__A1 (.I(_4433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4841__A2 (.I(_4433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8061__A2 (.I(_4434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7463__I (.I(_4434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7292__I (.I(_4434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4842__I (.I(_4434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8366__A3 (.I(_4435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8289__A2 (.I(_4435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7466__I (.I(_4435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4843__I (.I(_4435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8788__B2 (.I(_4436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8319__A2 (.I(_4436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7845__A1 (.I(_4436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4844__I (.I(_4436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7345__A1 (.I(_4437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7298__A2 (.I(_4437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5030__A1 (.I(_4437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4851__A3 (.I(_4437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5147__A2 (.I(_4438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5136__A1 (.I(_4438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5111__A1 (.I(_4438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4846__I (.I(_4438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7272__A2 (.I(_4439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6158__A1 (.I(_4439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5859__A1 (.I(_4439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4847__I (.I(_4439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7742__I (.I(_4440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7607__I (.I(_4440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6157__A1 (.I(_4440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4850__A1 (.I(_4440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7284__A1 (.I(_4441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7245__A1 (.I(_4441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4849__I (.I(_4441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8351__C (.I(_4443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7643__A1 (.I(_4443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4971__I (.I(_4443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4851__A4 (.I(_4443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4977__A1 (.I(_4444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4866__A2 (.I(_4444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6171__A2 (.I(_4445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6128__A2 (.I(_4445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4955__I (.I(_4445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4853__A2 (.I(_4445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5084__B1 (.I(_4446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4861__A1 (.I(_4446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7609__I (.I(_4447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7041__I (.I(_4447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5042__A2 (.I(_4447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4855__I (.I(_4447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8210__A2 (.I(_4448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8053__B (.I(_4448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7062__I (.I(_4448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4859__A1 (.I(_4448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6525__A1 (.I(_4449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6290__A1 (.I(_4449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5138__A1 (.I(_4449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4857__I (.I(_4449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7966__A1 (.I(_4450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6358__A1 (.I(_4450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6251__A3 (.I(_4450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4858__A1 (.I(_4450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8407__A1 (.I(\as2650.addr_buff[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8097__A1 (.I(\as2650.addr_buff[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7752__A3 (.I(\as2650.addr_buff[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7079__I (.I(\as2650.addr_buff[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8407__A2 (.I(\as2650.addr_buff[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8143__B2 (.I(\as2650.addr_buff[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7795__I (.I(\as2650.addr_buff[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7084__I (.I(\as2650.addr_buff[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4708__I (.I(\as2650.alu_op[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4576__A1 (.I(\as2650.alu_op[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4563__I (.I(\as2650.alu_op[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4576__A2 (.I(\as2650.alu_op[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4460__I (.I(\as2650.alu_op[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4634__I (.I(\as2650.alu_op[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4576__A3 (.I(\as2650.alu_op[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4564__A3 (.I(\as2650.alu_op[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5844__I (.I(\as2650.cycle[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5115__A2 (.I(\as2650.cycle[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5105__A1 (.I(\as2650.cycle[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4909__I (.I(\as2650.cycle[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4881__A1 (.I(\as2650.cycle[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4753__A2 (.I(\as2650.cycle[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4687__A2 (.I(\as2650.cycle[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5042__A1 (.I(\as2650.cycle[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4759__I (.I(\as2650.cycle[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4750__A2 (.I(\as2650.cycle[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4666__A2 (.I(\as2650.cycle[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4979__A2 (.I(\as2650.cycle[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4902__A1 (.I(\as2650.cycle[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4883__I (.I(\as2650.cycle[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4739__A2 (.I(\as2650.cycle[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5010__A1 (.I(\as2650.cycle[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4894__A2 (.I(\as2650.cycle[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4819__A1 (.I(\as2650.cycle[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4738__A2 (.I(\as2650.cycle[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5119__A2 (.I(\as2650.cycle[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4959__I (.I(\as2650.cycle[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4689__I (.I(\as2650.cycle[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5142__A1 (.I(\as2650.cycle[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4762__I (.I(\as2650.cycle[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4451__I (.I(\as2650.cycle[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4919__I (.I(\as2650.cycle[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4672__A2 (.I(\as2650.cycle[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5120__A2 (.I(\as2650.cycle[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5105__A2 (.I(\as2650.cycle[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4921__I (.I(\as2650.cycle[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4913__I (.I(\as2650.cycle[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5846__A1 (.I(\as2650.halted ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4715__A1 (.I(\as2650.halted ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4696__I (.I(\as2650.halted ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4649__I (.I(\as2650.halted ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5194__A1 (.I(\as2650.holding_reg[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5174__I (.I(\as2650.holding_reg[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7937__I1 (.I(\as2650.holding_reg[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5355__A1 (.I(\as2650.holding_reg[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5346__A1 (.I(\as2650.holding_reg[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5340__A1 (.I(\as2650.holding_reg[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7942__I1 (.I(\as2650.holding_reg[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5439__A1 (.I(\as2650.holding_reg[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5434__A1 (.I(\as2650.holding_reg[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5429__A1 (.I(\as2650.holding_reg[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7947__I1 (.I(\as2650.holding_reg[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5591__A1 (.I(\as2650.holding_reg[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5514__A1 (.I(\as2650.holding_reg[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5509__A1 (.I(\as2650.holding_reg[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7953__I1 (.I(\as2650.holding_reg[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5585__A1 (.I(\as2650.holding_reg[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5579__A1 (.I(\as2650.holding_reg[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5657__A1 (.I(\as2650.holding_reg[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5651__I (.I(\as2650.holding_reg[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7961__I1 (.I(\as2650.holding_reg[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5758__A1 (.I(\as2650.holding_reg[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5757__A1 (.I(\as2650.holding_reg[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5756__A1 (.I(\as2650.holding_reg[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7964__I1 (.I(\as2650.holding_reg[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5787__A1 (.I(\as2650.holding_reg[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5780__A1 (.I(\as2650.holding_reg[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5237__I (.I(\as2650.idx_ctrl[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5187__I (.I(\as2650.idx_ctrl[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5129__A2 (.I(\as2650.idx_ctrl[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5395__A1 (.I(\as2650.idx_ctrl[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5186__I (.I(\as2650.idx_ctrl[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5129__A1 (.I(\as2650.idx_ctrl[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4491__I (.I(\as2650.ins_reg[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4483__A2 (.I(\as2650.ins_reg[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4476__A2 (.I(\as2650.ins_reg[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4473__A2 (.I(\as2650.ins_reg[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4800__A2 (.I(\as2650.ins_reg[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4781__A2 (.I(\as2650.ins_reg[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4674__I (.I(\as2650.ins_reg[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4800__A1 (.I(\as2650.ins_reg[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4781__A1 (.I(\as2650.ins_reg[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4658__I (.I(\as2650.ins_reg[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4644__I (.I(\as2650.ins_reg[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8873__A1 (.I(\as2650.overflow ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8540__A1 (.I(\as2650.overflow ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6381__A1 (.I(\as2650.overflow ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7791__A1 (.I(\as2650.pc[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6031__I (.I(\as2650.pc[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7836__A1 (.I(\as2650.pc[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7820__I (.I(\as2650.pc[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6042__I (.I(\as2650.pc[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8456__A1 (.I(\as2650.pc[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8451__A1 (.I(\as2650.pc[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6057__I (.I(\as2650.pc[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7377__A1 (.I(\as2650.pc[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7330__A1 (.I(\as2650.pc[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7323__I (.I(\as2650.pc[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5886__I (.I(\as2650.pc[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8126__A1 (.I(\as2650.pc[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7405__I (.I(\as2650.pc[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7375__A1 (.I(\as2650.pc[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5892__I (.I(\as2650.pc[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7453__I (.I(\as2650.pc[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7444__A1 (.I(\as2650.pc[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5897__I (.I(\as2650.pc[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8308__A2 (.I(\as2650.pc[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7686__A1 (.I(\as2650.pc[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7626__I (.I(\as2650.pc[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5932__I (.I(\as2650.pc[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8357__A1 (.I(\as2650.pc[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7766__A1 (.I(\as2650.pc[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7714__I (.I(\as2650.pc[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6012__I (.I(\as2650.pc[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8888__B (.I(\as2650.psl[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8522__A1 (.I(\as2650.psl[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6377__A1 (.I(\as2650.psl[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6269__A1 (.I(\as2650.psl[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5209__A1 (.I(\as2650.psl[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5199__I (.I(\as2650.psl[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6540__S (.I(\as2650.psl[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4494__I (.I(\as2650.psl[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4467__I (.I(\as2650.psl[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8864__A1 (.I(\as2650.psl[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8587__A1 (.I(\as2650.psl[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6381__B2 (.I(\as2650.psl[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6373__A1 (.I(\as2650.psl[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6352__I (.I(\as2650.psl[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4629__A1 (.I(\as2650.psl[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7184__A2 (.I(\as2650.psu[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5302__A2 (.I(\as2650.psu[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5298__I (.I(\as2650.psu[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5291__I (.I(\as2650.psu[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6387__B2 (.I(\as2650.psu[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5964__I (.I(\as2650.psu[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5497__A1 (.I(\as2650.psu[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5310__I (.I(\as2650.psu[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8900__B (.I(\as2650.psu[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8556__A1 (.I(\as2650.psu[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6386__B2 (.I(\as2650.psu[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8897__B (.I(\as2650.psu[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8574__A1 (.I(\as2650.psu[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6385__I (.I(\as2650.psu[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8586__A1 (.I(\as2650.psu[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6389__A1 (.I(\as2650.psu[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6149__A1 (.I(\as2650.psu[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6103__I (.I(\as2650.psu[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8616__A1 (.I(\as2650.psu[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7969__I (.I(\as2650.psu[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6387__C1 (.I(\as2650.psu[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6633__A1 (.I(\as2650.r0[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4565__I (.I(\as2650.r0[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6668__A1 (.I(\as2650.r0[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6631__A1 (.I(\as2650.r0[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4555__I (.I(\as2650.r0[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6707__A1 (.I(\as2650.r0[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6672__A1 (.I(\as2650.r0[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6632__A1 (.I(\as2650.r0[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4544__I (.I(\as2650.r0[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6764__A1 (.I(\as2650.r0[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6671__A1 (.I(\as2650.r0[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4533__I (.I(\as2650.r0[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6815__B2 (.I(\as2650.r0[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6767__A1 (.I(\as2650.r0[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4523__I (.I(\as2650.r0[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6813__A1 (.I(\as2650.r0[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6651__I (.I(\as2650.r0[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4511__I (.I(\as2650.r0[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6636__A1 (.I(\as2650.r0[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4504__I (.I(\as2650.r0[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6665__A1 (.I(\as2650.r0[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4481__I (.I(\as2650.r0[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6551__I0 (.I(\as2650.r123[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6007__A1 (.I(\as2650.r123[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5104__I (.I(\as2650.r123[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4568__I1 (.I(\as2650.r123[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6554__I0 (.I(\as2650.r123[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6018__A1 (.I(\as2650.r123[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5338__I (.I(\as2650.r123[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4551__I1 (.I(\as2650.r123[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6572__I0 (.I(\as2650.r123[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6027__A1 (.I(\as2650.r123[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5428__I (.I(\as2650.r123[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4546__I1 (.I(\as2650.r123[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6557__I0 (.I(\as2650.r123[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6038__A1 (.I(\as2650.r123[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5505__I (.I(\as2650.r123[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4537__I1 (.I(\as2650.r123[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6543__I0 (.I(\as2650.r123[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6045__A1 (.I(\as2650.r123[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5576__I (.I(\as2650.r123[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4528__I1 (.I(\as2650.r123[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6540__I0 (.I(\as2650.r123[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6053__A1 (.I(\as2650.r123[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5649__I (.I(\as2650.r123[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4519__I1 (.I(\as2650.r123[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6061__A1 (.I(\as2650.r123[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5715__I (.I(\as2650.r123[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4495__I0 (.I(\as2650.r123[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8722__A1 (.I(\as2650.r123[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4528__I0 (.I(\as2650.r123[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8728__B2 (.I(\as2650.r123[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4519__I0 (.I(\as2650.r123[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8730__B2 (.I(\as2650.r123[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4490__I (.I(\as2650.r123[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8732__B2 (.I(\as2650.r123[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4471__I0 (.I(\as2650.r123[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7140__A1 (.I(\as2650.r123_2[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6551__I1 (.I(\as2650.r123_2[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5999__A1 (.I(\as2650.r123_2[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4568__I3 (.I(\as2650.r123_2[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7150__A1 (.I(\as2650.r123_2[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6554__I1 (.I(\as2650.r123_2[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6016__A1 (.I(\as2650.r123_2[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4551__I3 (.I(\as2650.r123_2[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7156__A1 (.I(\as2650.r123_2[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6572__I1 (.I(\as2650.r123_2[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6025__A1 (.I(\as2650.r123_2[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4546__I3 (.I(\as2650.r123_2[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7161__A1 (.I(\as2650.r123_2[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6557__I1 (.I(\as2650.r123_2[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6036__A1 (.I(\as2650.r123_2[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4537__I3 (.I(\as2650.r123_2[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7167__A1 (.I(\as2650.r123_2[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6543__I1 (.I(\as2650.r123_2[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6043__A1 (.I(\as2650.r123_2[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4528__I3 (.I(\as2650.r123_2[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7172__A1 (.I(\as2650.r123_2[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6540__I1 (.I(\as2650.r123_2[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6051__A1 (.I(\as2650.r123_2[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4519__I3 (.I(\as2650.r123_2[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7174__A1 (.I(\as2650.r123_2[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6059__A1 (.I(\as2650.r123_2[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4495__I1 (.I(\as2650.r123_2[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7004__B2 (.I(\as2650.r123_2[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4568__I2 (.I(\as2650.r123_2[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7011__A1 (.I(\as2650.r123_2[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4551__I2 (.I(\as2650.r123_2[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7026__A1 (.I(\as2650.r123_2[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4519__I2 (.I(\as2650.r123_2[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7030__A1 (.I(\as2650.r123_2[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4489__A2 (.I(\as2650.r123_2[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7033__A1 (.I(\as2650.r123_2[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4471__I2 (.I(\as2650.r123_2[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6828__A1 (.I(\as2650.r123_2[2][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4541__I1 (.I(\as2650.r123_2[2][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6447__A1 (.I(\as2650.stack[0][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5499__B2 (.I(\as2650.stack[0][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6455__A1 (.I(\as2650.stack[0][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5722__B2 (.I(\as2650.stack[0][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6029__A1 (.I(\as2650.stack[1][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5499__A1 (.I(\as2650.stack[1][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6063__A1 (.I(\as2650.stack[1][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5722__A1 (.I(\as2650.stack[1][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8278__A1 (.I(\as2650.stack[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5986__A1 (.I(\as2650.stack[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8014__B2 (.I(\as2650.stack[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5942__A1 (.I(\as2650.stack[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8074__B2 (.I(\as2650.stack[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5944__A1 (.I(\as2650.stack[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8117__B2 (.I(\as2650.stack[2][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5946__A1 (.I(\as2650.stack[2][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8261__B2 (.I(\as2650.stack[2][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5956__A1 (.I(\as2650.stack[2][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8277__B2 (.I(\as2650.stack[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5958__A1 (.I(\as2650.stack[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8199__A1 (.I(\as2650.stack[3][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5921__A1 (.I(\as2650.stack[3][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8261__A1 (.I(\as2650.stack[3][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5930__A1 (.I(\as2650.stack[3][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8277__A1 (.I(\as2650.stack[3][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5937__A1 (.I(\as2650.stack[3][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8763__A1 (.I(\as2650.stack[4][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8022__A1 (.I(\as2650.stack[4][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8767__A1 (.I(\as2650.stack[4][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8115__B2 (.I(\as2650.stack[4][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8773__A1 (.I(\as2650.stack[4][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8185__B2 (.I(\as2650.stack[4][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8779__A1 (.I(\as2650.stack[4][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8281__B2 (.I(\as2650.stack[4][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8185__A1 (.I(\as2650.stack[5][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6989__A1 (.I(\as2650.stack[5][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8263__A1 (.I(\as2650.stack[5][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6995__A1 (.I(\as2650.stack[5][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8279__A1 (.I(\as2650.stack[5][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6998__A1 (.I(\as2650.stack[5][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8666__A1 (.I(\as2650.stack[6][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8020__B2 (.I(\as2650.stack[6][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8668__A1 (.I(\as2650.stack[6][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8072__B2 (.I(\as2650.stack[6][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8676__A1 (.I(\as2650.stack[6][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8184__B2 (.I(\as2650.stack[6][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8628__A1 (.I(\as2650.stack[7][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8072__A1 (.I(\as2650.stack[7][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1_I (.I(io_in[10]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input2_I (.I(io_in[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input3_I (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input4_I (.I(io_in[13]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input5_I (.I(io_in[33]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input6_I (.I(io_in[34]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input7_I (.I(io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input8_I (.I(io_in[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input9_I (.I(io_in[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input10_I (.I(io_in[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input11_I (.I(io_in[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9008__CLK (.I(clknet_leaf_1_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9093__CLK (.I(clknet_leaf_1_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9096__CLK (.I(clknet_leaf_1_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8987__CLK (.I(clknet_leaf_1_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_0_wb_clk_i_I (.I(wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6145__I (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5686__I (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6317__I (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5736__I (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7325__I (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5811__I (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4966__I (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4820__I (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7972__B (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4715__A2 (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4665__I (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4650__I (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4750__A1 (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4669__I (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4666__A1 (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8051__A1 (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7363__A2 (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7329__A2 (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5265__I (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7330__A2 (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5375__I (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7375__A2 (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5473__I (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7480__I (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6371__I (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5545__I (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7602__A2 (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7517__A2 (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7479__A2 (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5613__I (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output12_I (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output15_I (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output16_I (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output17_I (.I(net17));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output18_I (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output20_I (.I(net20));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6215__A1 (.I(net20));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output21_I (.I(net21));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6219__A1 (.I(net21));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output22_I (.I(net22));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6224__A1 (.I(net22));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output25_I (.I(net25));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7214__A1 (.I(net25));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout52_I (.I(net26));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output26_I (.I(net26));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output27_I (.I(net27));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7870__C2 (.I(net27));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5087__I (.I(net27));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output28_I (.I(net28));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8893__B (.I(net28));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8602__I (.I(net28));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6389__B2 (.I(net28));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output29_I (.I(net29));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7439__A3 (.I(net29));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7280__I (.I(net29));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output30_I (.I(net30));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7439__A2 (.I(net30));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7373__A1 (.I(net30));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7333__I (.I(net30));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output31_I (.I(net31));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7439__A1 (.I(net31));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7372__I (.I(net31));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output33_I (.I(net33));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7555__A1 (.I(net33));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7484__I (.I(net33));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output34_I (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7636__A2 (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7595__A1 (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7554__I (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output35_I (.I(net35));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7636__A1 (.I(net35));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7578__I (.I(net35));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout54_I (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output36_I (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output37_I (.I(net37));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7760__A2 (.I(net37));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7728__A1 (.I(net37));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7679__I (.I(net37));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output38_I (.I(net38));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7760__A1 (.I(net38));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7727__I (.I(net38));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output39_I (.I(net39));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7801__I (.I(net39));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7759__I (.I(net39));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output40_I (.I(net40));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7828__A1 (.I(net40));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7800__I (.I(net40));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout53_I (.I(net41));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output41_I (.I(net41));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output42_I (.I(net42));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6185__A1 (.I(net42));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9240__I (.I(net48));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9239__I (.I(net48));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9238__I (.I(net48));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7904__A1 (.I(net52));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7900__A1 (.I(net52));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7899__A1 (.I(net52));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7897__A1 (.I(net52));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7851__A1 (.I(net53));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7844__A1 (.I(net53));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7842__A1 (.I(net53));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7829__A1 (.I(net53));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7666__A1 (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7640__A1 (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7637__A1 (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7632__I (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7477__A1 (.I(net55));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7468__A1 (.I(net55));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7454__I (.I(net55));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7440__A1 (.I(net55));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9157__CLK (.I(clknet_leaf_3_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8986__CLK (.I(clknet_leaf_3_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9024__CLK (.I(clknet_leaf_5_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9022__CLK (.I(clknet_leaf_5_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9021__CLK (.I(clknet_leaf_5_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9170__CLK (.I(clknet_leaf_5_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9091__CLK (.I(clknet_leaf_9_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9033__CLK (.I(clknet_leaf_9_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9090__CLK (.I(clknet_leaf_9_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9034__CLK (.I(clknet_leaf_9_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8988__CLK (.I(clknet_leaf_9_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8989__CLK (.I(clknet_leaf_9_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9043__CLK (.I(clknet_leaf_15_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8970__CLK (.I(clknet_leaf_15_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8969__CLK (.I(clknet_leaf_15_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8971__CLK (.I(clknet_leaf_15_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8972__CLK (.I(clknet_leaf_15_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8967__CLK (.I(clknet_leaf_15_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8968__CLK (.I(clknet_leaf_15_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9102__CLK (.I(clknet_leaf_15_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9088__CLK (.I(clknet_leaf_16_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8974__CLK (.I(clknet_leaf_16_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8973__CLK (.I(clknet_leaf_16_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9089__CLK (.I(clknet_leaf_17_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9073__CLK (.I(clknet_leaf_17_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9072__CLK (.I(clknet_leaf_17_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9082__CLK (.I(clknet_leaf_22_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9083__CLK (.I(clknet_leaf_22_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9078__CLK (.I(clknet_leaf_22_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9081__CLK (.I(clknet_leaf_22_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9112__CLK (.I(clknet_leaf_27_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9111__CLK (.I(clknet_leaf_27_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9109__CLK (.I(clknet_leaf_27_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9104__CLK (.I(clknet_leaf_27_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9049__CLK (.I(clknet_leaf_29_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9114__CLK (.I(clknet_leaf_29_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9016__CLK (.I(clknet_leaf_30_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9017__CLK (.I(clknet_leaf_30_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9131__CLK (.I(clknet_leaf_30_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9145__CLK (.I(clknet_leaf_30_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9144__CLK (.I(clknet_leaf_30_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8932__CLK (.I(clknet_leaf_31_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8933__CLK (.I(clknet_leaf_31_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8934__CLK (.I(clknet_leaf_31_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9175__CLK (.I(clknet_leaf_31_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9176__CLK (.I(clknet_leaf_31_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9178__CLK (.I(clknet_leaf_31_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9177__CLK (.I(clknet_leaf_31_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9018__CLK (.I(clknet_leaf_31_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9019__CLK (.I(clknet_leaf_31_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8931__CLK (.I(clknet_leaf_32_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8923__CLK (.I(clknet_leaf_32_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8926__CLK (.I(clknet_leaf_32_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8924__CLK (.I(clknet_leaf_32_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8925__CLK (.I(clknet_leaf_32_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9132__CLK (.I(clknet_leaf_33_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9130__CLK (.I(clknet_leaf_33_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9129__CLK (.I(clknet_leaf_33_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8954__CLK (.I(clknet_leaf_33_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9014__CLK (.I(clknet_leaf_34_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9012__CLK (.I(clknet_leaf_34_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9125__CLK (.I(clknet_leaf_34_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9147__CLK (.I(clknet_leaf_34_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9146__CLK (.I(clknet_leaf_34_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9128__CLK (.I(clknet_leaf_34_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9171__CLK (.I(clknet_leaf_36_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9174__CLK (.I(clknet_leaf_36_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9173__CLK (.I(clknet_leaf_36_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9172__CLK (.I(clknet_leaf_36_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8927__CLK (.I(clknet_leaf_36_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8930__CLK (.I(clknet_leaf_36_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9142__CLK (.I(clknet_leaf_37_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9143__CLK (.I(clknet_leaf_37_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9140__CLK (.I(clknet_leaf_37_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9141__CLK (.I(clknet_leaf_37_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9100__CLK (.I(clknet_leaf_37_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9115__CLK (.I(clknet_leaf_38_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9126__CLK (.I(clknet_leaf_38_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9127__CLK (.I(clknet_leaf_38_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9182__CLK (.I(clknet_leaf_41_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9183__CLK (.I(clknet_leaf_41_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8928__CLK (.I(clknet_leaf_41_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8929__CLK (.I(clknet_leaf_41_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9189__CLK (.I(clknet_leaf_43_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9190__CLK (.I(clknet_leaf_43_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8966__CLK (.I(clknet_leaf_43_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9154__CLK (.I(clknet_leaf_44_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9056__CLK (.I(clknet_leaf_44_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9139__CLK (.I(clknet_leaf_44_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9138__CLK (.I(clknet_leaf_44_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9003__CLK (.I(clknet_leaf_44_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9188__CLK (.I(clknet_leaf_44_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9186__CLK (.I(clknet_leaf_44_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9181__CLK (.I(clknet_leaf_45_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9153__CLK (.I(clknet_leaf_45_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9191__CLK (.I(clknet_leaf_45_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9192__CLK (.I(clknet_leaf_45_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9055__CLK (.I(clknet_leaf_45_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9001__CLK (.I(clknet_leaf_46_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9133__CLK (.I(clknet_leaf_46_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9148__CLK (.I(clknet_leaf_46_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9050__CLK (.I(clknet_leaf_46_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9054__CLK (.I(clknet_leaf_46_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9152__CLK (.I(clknet_leaf_46_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8949__CLK (.I(clknet_leaf_48_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8948__CLK (.I(clknet_leaf_48_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8980__CLK (.I(clknet_leaf_48_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9070__CLK (.I(clknet_leaf_48_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9071__CLK (.I(clknet_leaf_48_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9002__CLK (.I(clknet_leaf_48_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9065__CLK (.I(clknet_leaf_49_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8996__CLK (.I(clknet_leaf_49_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8979__CLK (.I(clknet_leaf_50_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8947__CLK (.I(clknet_leaf_50_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8990__CLK (.I(clknet_leaf_50_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8994__CLK (.I(clknet_leaf_50_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8943__CLK (.I(clknet_leaf_50_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9069__CLK (.I(clknet_leaf_50_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8977__CLK (.I(clknet_leaf_51_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8991__CLK (.I(clknet_leaf_51_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8944__CLK (.I(clknet_leaf_51_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8976__CLK (.I(clknet_leaf_51_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9066__CLK (.I(clknet_leaf_51_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8978__CLK (.I(clknet_leaf_51_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8952__CLK (.I(clknet_leaf_54_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8950__CLK (.I(clknet_leaf_54_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8953__CLK (.I(clknet_leaf_54_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8951__CLK (.I(clknet_leaf_54_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9051__CLK (.I(clknet_leaf_54_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8922__CLK (.I(clknet_leaf_54_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8956__CLK (.I(clknet_leaf_57_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8957__CLK (.I(clknet_leaf_57_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8955__CLK (.I(clknet_leaf_57_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8935__CLK (.I(clknet_leaf_57_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8993__CLK (.I(clknet_leaf_59_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8992__CLK (.I(clknet_leaf_59_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8946__CLK (.I(clknet_leaf_59_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8945__CLK (.I(clknet_leaf_59_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9068__CLK (.I(clknet_leaf_59_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9187__CLK (.I(clknet_leaf_67_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8995__CLK (.I(clknet_leaf_67_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8914__CLK (.I(clknet_leaf_68_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8911__CLK (.I(clknet_leaf_68_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8917__CLK (.I(clknet_leaf_68_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8912__CLK (.I(clknet_leaf_68_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8913__CLK (.I(clknet_leaf_68_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8915__CLK (.I(clknet_leaf_68_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8916__CLK (.I(clknet_leaf_68_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9062__CLK (.I(clknet_leaf_70_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9059__CLK (.I(clknet_leaf_70_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9060__CLK (.I(clknet_leaf_70_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9063__CLK (.I(clknet_leaf_70_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9058__CLK (.I(clknet_leaf_70_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9064__CLK (.I(clknet_leaf_70_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9057__CLK (.I(clknet_leaf_70_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9061__CLK (.I(clknet_leaf_70_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9160__CLK (.I(clknet_leaf_71_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9155__CLK (.I(clknet_leaf_71_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9162__CLK (.I(clknet_leaf_71_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9025__CLK (.I(clknet_leaf_71_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9004__CLK (.I(clknet_leaf_77_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9163__CLK (.I(clknet_leaf_77_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9011__CLK (.I(clknet_leaf_77_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9010__CLK (.I(clknet_leaf_77_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9123__CLK (.I(clknet_leaf_82_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9097__CLK (.I(clknet_leaf_82_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9094__CLK (.I(clknet_leaf_82_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9184__CLK (.I(clknet_leaf_82_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9098__CLK (.I(clknet_leaf_82_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9099__CLK (.I(clknet_leaf_82_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_7__f_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_6__f_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_5__f_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_4__f_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_3__f_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_2__f_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_1__f_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_0__f_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_82_wb_clk_i_I (.I(clknet_3_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_81_wb_clk_i_I (.I(clknet_3_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_80_wb_clk_i_I (.I(clknet_3_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_79_wb_clk_i_I (.I(clknet_3_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_78_wb_clk_i_I (.I(clknet_3_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_77_wb_clk_i_I (.I(clknet_3_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_76_wb_clk_i_I (.I(clknet_3_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_4_wb_clk_i_I (.I(clknet_3_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_2_wb_clk_i_I (.I(clknet_3_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9095__CLK (.I(clknet_3_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_75_wb_clk_i_I (.I(clknet_3_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_74_wb_clk_i_I (.I(clknet_3_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_73_wb_clk_i_I (.I(clknet_3_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8918__CLK (.I(clknet_3_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_71_wb_clk_i_I (.I(clknet_3_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_70_wb_clk_i_I (.I(clknet_3_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_69_wb_clk_i_I (.I(clknet_3_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8982__CLK (.I(clknet_3_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_7_wb_clk_i_I (.I(clknet_3_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_6_wb_clk_i_I (.I(clknet_3_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_5_wb_clk_i_I (.I(clknet_3_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_16_wb_clk_i_I (.I(clknet_3_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_15_wb_clk_i_I (.I(clknet_3_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_14_wb_clk_i_I (.I(clknet_3_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_13_wb_clk_i_I (.I(clknet_3_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9047__CLK (.I(clknet_3_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9040__CLK (.I(clknet_3_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9180__CLK (.I(clknet_3_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_9_wb_clk_i_I (.I(clknet_3_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_1_wb_clk_i_I (.I(clknet_3_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_21_wb_clk_i_I (.I(clknet_3_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_20_wb_clk_i_I (.I(clknet_3_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_opt_2_0_wb_clk_i_I (.I(clknet_3_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_18_wb_clk_i_I (.I(clknet_3_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_17_wb_clk_i_I (.I(clknet_3_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_opt_1_0_wb_clk_i_I (.I(clknet_3_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_68_wb_clk_i_I (.I(clknet_3_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_67_wb_clk_i_I (.I(clknet_3_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_59_wb_clk_i_I (.I(clknet_3_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_51_wb_clk_i_I (.I(clknet_3_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_50_wb_clk_i_I (.I(clknet_3_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_49_wb_clk_i_I (.I(clknet_3_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_48_wb_clk_i_I (.I(clknet_3_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_47_wb_clk_i_I (.I(clknet_3_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_46_wb_clk_i_I (.I(clknet_3_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_45_wb_clk_i_I (.I(clknet_3_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_44_wb_clk_i_I (.I(clknet_3_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_43_wb_clk_i_I (.I(clknet_3_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_66_wb_clk_i_I (.I(clknet_3_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8962__CLK (.I(clknet_3_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8961__CLK (.I(clknet_3_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_63_wb_clk_i_I (.I(clknet_3_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8963__CLK (.I(clknet_3_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_61_wb_clk_i_I (.I(clknet_3_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_60_wb_clk_i_I (.I(clknet_3_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_40_wb_clk_i_I (.I(clknet_3_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9116__CLK (.I(clknet_3_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_38_wb_clk_i_I (.I(clknet_3_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_37_wb_clk_i_I (.I(clknet_3_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_29_wb_clk_i_I (.I(clknet_3_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9113__CLK (.I(clknet_3_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_27_wb_clk_i_I (.I(clknet_3_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9103__CLK (.I(clknet_3_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_25_wb_clk_i_I (.I(clknet_3_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_24_wb_clk_i_I (.I(clknet_3_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_opt_4_0_wb_clk_i_I (.I(clknet_3_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_opt_3_0_wb_clk_i_I (.I(clknet_3_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_58_wb_clk_i_I (.I(clknet_3_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_57_wb_clk_i_I (.I(clknet_3_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_56_wb_clk_i_I (.I(clknet_3_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_55_wb_clk_i_I (.I(clknet_3_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_54_wb_clk_i_I (.I(clknet_3_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_53_wb_clk_i_I (.I(clknet_3_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_52_wb_clk_i_I (.I(clknet_3_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9185__CLK (.I(clknet_3_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_41_wb_clk_i_I (.I(clknet_3_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_36_wb_clk_i_I (.I(clknet_3_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_35_wb_clk_i_I (.I(clknet_3_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_34_wb_clk_i_I (.I(clknet_3_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_33_wb_clk_i_I (.I(clknet_3_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_32_wb_clk_i_I (.I(clknet_3_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_31_wb_clk_i_I (.I(clknet_3_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_30_wb_clk_i_I (.I(clknet_3_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_3_wb_clk_i_I (.I(clknet_opt_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_19_wb_clk_i_I (.I(clknet_opt_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_22_wb_clk_i_I (.I(clknet_opt_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_23_wb_clk_i_I (.I(clknet_opt_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_9_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_11_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_15_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_17_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_30_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_30_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_33_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_33_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_33_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_33_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_35_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_35_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_37_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_39_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_43_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_43_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_45_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_45_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_47_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_47_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_47_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_47_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_48_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_48_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_49_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_55_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_55_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_57_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_57_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_59_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_59_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_59_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_59_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_59_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_61_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_61_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_63_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_63_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_63_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_63_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_63_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_63_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_63_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_63_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_63_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_65_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_69_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_69_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_69_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_70_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_70_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_70_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_70_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_71_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_71_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_71_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_71_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_71_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_72_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_72_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_72_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_73_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_73_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_73_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_75_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_75_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_75_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_75_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_75_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_77_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_77_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_79_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_79_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_79_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_79_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_79_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_79_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_81_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_81_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_81_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_89_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_89_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_89_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_89_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_89_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_89_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_91_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_91_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_91_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_91_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_93_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_93_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_93_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_93_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_95_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_95_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_95_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_95_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_95_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_95_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_95_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_95_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_97_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_97_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_97_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_97_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_97_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_99_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_99_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_99_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_101_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_101_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_101_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_101_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_101_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_103_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_103_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_103_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_103_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_103_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_103_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_105_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_105_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_105_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_105_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_105_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_105_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_107_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_107_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_107_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_107_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_109_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_109_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_109_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_111_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_111_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_111_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_113_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_113_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_113_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_113_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_113_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_113_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_115_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_117_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_117_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_117_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_117_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_117_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_117_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_117_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_117_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_119_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_119_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_119_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_121_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_121_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_121_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_121_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_121_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_121_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_123_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_123_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_123_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_127_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_127_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_127_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_127_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_127_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_127_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_129_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_131_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_131_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_131_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_131_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_133_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_135_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_135_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_135_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_135_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_135_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_135_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_135_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_135_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_137_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_139_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_139_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_139_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_139_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_140_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_140_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_140_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_140_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_140_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_141_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_141_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_143_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_143_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_143_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1577 ();
 assign io_oeb[0] = net86;
 assign io_oeb[13] = net91;
 assign io_oeb[14] = net56;
 assign io_oeb[15] = net57;
 assign io_oeb[16] = net58;
 assign io_oeb[17] = net59;
 assign io_oeb[18] = net60;
 assign io_oeb[19] = net61;
 assign io_oeb[1] = net87;
 assign io_oeb[20] = net62;
 assign io_oeb[21] = net63;
 assign io_oeb[22] = net64;
 assign io_oeb[23] = net65;
 assign io_oeb[24] = net66;
 assign io_oeb[25] = net67;
 assign io_oeb[26] = net68;
 assign io_oeb[27] = net69;
 assign io_oeb[28] = net70;
 assign io_oeb[29] = net71;
 assign io_oeb[2] = net88;
 assign io_oeb[30] = net72;
 assign io_oeb[31] = net73;
 assign io_oeb[32] = net74;
 assign io_oeb[33] = net92;
 assign io_oeb[34] = net93;
 assign io_oeb[35] = net94;
 assign io_oeb[36] = net95;
 assign io_oeb[37] = net96;
 assign io_oeb[3] = net89;
 assign io_oeb[4] = net90;
 assign io_out[0] = net75;
 assign io_out[13] = net80;
 assign io_out[1] = net76;
 assign io_out[2] = net77;
 assign io_out[33] = net81;
 assign io_out[34] = net82;
 assign io_out[35] = net83;
 assign io_out[36] = net84;
 assign io_out[37] = net85;
 assign io_out[3] = net78;
 assign io_out[4] = net79;
endmodule

