magic
tech gf180mcuD
magscale 1 5
timestamp 1700266336
<< obsm1 >>
rect 672 1538 41776 40798
<< metal2 >>
rect 4144 42100 4200 42500
rect 12656 42100 12712 42500
rect 21168 42100 21224 42500
rect 29680 42100 29736 42500
rect 38192 42100 38248 42500
rect 2352 0 2408 400
rect 7056 0 7112 400
rect 11760 0 11816 400
rect 16464 0 16520 400
rect 21168 0 21224 400
rect 25872 0 25928 400
rect 30576 0 30632 400
rect 35280 0 35336 400
rect 39984 0 40040 400
<< obsm2 >>
rect 574 42070 4114 42100
rect 4230 42070 12626 42100
rect 12742 42070 21138 42100
rect 21254 42070 29650 42100
rect 29766 42070 38162 42100
rect 38278 42070 41594 42100
rect 574 430 41594 42070
rect 574 400 2322 430
rect 2438 400 7026 430
rect 7142 400 11730 430
rect 11846 400 16434 430
rect 16550 400 21138 430
rect 21254 400 25842 430
rect 25958 400 30546 430
rect 30662 400 35250 430
rect 35366 400 39954 430
rect 40070 400 41594 430
<< metal3 >>
rect 0 40880 400 40936
rect 42100 39648 42500 39704
rect 0 37856 400 37912
rect 0 34832 400 34888
rect 42100 34384 42500 34440
rect 0 31808 400 31864
rect 42100 29120 42500 29176
rect 0 28784 400 28840
rect 0 25760 400 25816
rect 42100 23856 42500 23912
rect 0 22736 400 22792
rect 0 19712 400 19768
rect 42100 18592 42500 18648
rect 0 16688 400 16744
rect 0 13664 400 13720
rect 42100 13328 42500 13384
rect 0 10640 400 10696
rect 42100 8064 42500 8120
rect 0 7616 400 7672
rect 0 4592 400 4648
rect 42100 2800 42500 2856
rect 0 1568 400 1624
<< obsm3 >>
rect 430 40850 42100 40922
rect 400 39734 42100 40850
rect 400 39618 42070 39734
rect 400 37942 42100 39618
rect 430 37826 42100 37942
rect 400 34918 42100 37826
rect 430 34802 42100 34918
rect 400 34470 42100 34802
rect 400 34354 42070 34470
rect 400 31894 42100 34354
rect 430 31778 42100 31894
rect 400 29206 42100 31778
rect 400 29090 42070 29206
rect 400 28870 42100 29090
rect 430 28754 42100 28870
rect 400 25846 42100 28754
rect 430 25730 42100 25846
rect 400 23942 42100 25730
rect 400 23826 42070 23942
rect 400 22822 42100 23826
rect 430 22706 42100 22822
rect 400 19798 42100 22706
rect 430 19682 42100 19798
rect 400 18678 42100 19682
rect 400 18562 42070 18678
rect 400 16774 42100 18562
rect 430 16658 42100 16774
rect 400 13750 42100 16658
rect 430 13634 42100 13750
rect 400 13414 42100 13634
rect 400 13298 42070 13414
rect 400 10726 42100 13298
rect 430 10610 42100 10726
rect 400 8150 42100 10610
rect 400 8034 42070 8150
rect 400 7702 42100 8034
rect 430 7586 42100 7702
rect 400 4678 42100 7586
rect 430 4562 42100 4678
rect 400 2886 42100 4562
rect 400 2770 42070 2886
rect 400 1654 42100 2770
rect 430 1554 42100 1654
<< metal4 >>
rect 2224 1538 2384 40798
rect 9904 1538 10064 40798
rect 17584 1538 17744 40798
rect 25264 1538 25424 40798
rect 32944 1538 33104 40798
rect 40624 1538 40784 40798
<< obsm4 >>
rect 2422 2977 9874 38519
rect 10094 2977 17554 38519
rect 17774 2977 25234 38519
rect 25454 2977 32914 38519
rect 33134 2977 39074 38519
<< labels >>
rlabel metal3 s 0 1568 400 1624 6 addr[0]
port 1 nsew signal input
rlabel metal3 s 0 4592 400 4648 6 addr[1]
port 2 nsew signal input
rlabel metal3 s 0 7616 400 7672 6 addr[2]
port 3 nsew signal input
rlabel metal3 s 0 10640 400 10696 6 addr[3]
port 4 nsew signal input
rlabel metal3 s 0 13664 400 13720 6 addr[4]
port 5 nsew signal input
rlabel metal3 s 0 16688 400 16744 6 addr[5]
port 6 nsew signal input
rlabel metal2 s 2352 0 2408 400 6 bus_cyc
port 7 nsew signal input
rlabel metal2 s 7056 0 7112 400 6 bus_we
port 8 nsew signal input
rlabel metal3 s 0 19712 400 19768 6 data_in[0]
port 9 nsew signal input
rlabel metal3 s 0 22736 400 22792 6 data_in[1]
port 10 nsew signal input
rlabel metal3 s 0 25760 400 25816 6 data_in[2]
port 11 nsew signal input
rlabel metal3 s 0 28784 400 28840 6 data_in[3]
port 12 nsew signal input
rlabel metal3 s 0 31808 400 31864 6 data_in[4]
port 13 nsew signal input
rlabel metal3 s 0 34832 400 34888 6 data_in[5]
port 14 nsew signal input
rlabel metal3 s 0 37856 400 37912 6 data_in[6]
port 15 nsew signal input
rlabel metal3 s 0 40880 400 40936 6 data_in[7]
port 16 nsew signal input
rlabel metal3 s 42100 2800 42500 2856 6 data_out[0]
port 17 nsew signal output
rlabel metal3 s 42100 8064 42500 8120 6 data_out[1]
port 18 nsew signal output
rlabel metal3 s 42100 13328 42500 13384 6 data_out[2]
port 19 nsew signal output
rlabel metal3 s 42100 18592 42500 18648 6 data_out[3]
port 20 nsew signal output
rlabel metal3 s 42100 23856 42500 23912 6 data_out[4]
port 21 nsew signal output
rlabel metal3 s 42100 29120 42500 29176 6 data_out[5]
port 22 nsew signal output
rlabel metal3 s 42100 34384 42500 34440 6 data_out[6]
port 23 nsew signal output
rlabel metal3 s 42100 39648 42500 39704 6 data_out[7]
port 24 nsew signal output
rlabel metal2 s 11760 0 11816 400 6 irq1
port 25 nsew signal output
rlabel metal2 s 16464 0 16520 400 6 irq2
port 26 nsew signal output
rlabel metal2 s 21168 0 21224 400 6 irq5
port 27 nsew signal output
rlabel metal2 s 21168 42100 21224 42500 6 pwm0
port 28 nsew signal output
rlabel metal2 s 29680 42100 29736 42500 6 pwm1
port 29 nsew signal output
rlabel metal2 s 38192 42100 38248 42500 6 pwm2
port 30 nsew signal output
rlabel metal2 s 30576 0 30632 400 6 rst
port 31 nsew signal input
rlabel metal2 s 35280 0 35336 400 6 tmr0_clk
port 32 nsew signal input
rlabel metal2 s 4144 42100 4200 42500 6 tmr0_o
port 33 nsew signal output
rlabel metal2 s 39984 0 40040 400 6 tmr1_clk
port 34 nsew signal input
rlabel metal2 s 12656 42100 12712 42500 6 tmr1_o
port 35 nsew signal output
rlabel metal4 s 2224 1538 2384 40798 6 vdd
port 36 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 40798 6 vdd
port 36 nsew power bidirectional
rlabel metal4 s 32944 1538 33104 40798 6 vdd
port 36 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 40798 6 vss
port 37 nsew ground bidirectional
rlabel metal4 s 25264 1538 25424 40798 6 vss
port 37 nsew ground bidirectional
rlabel metal4 s 40624 1538 40784 40798 6 vss
port 37 nsew ground bidirectional
rlabel metal2 s 25872 0 25928 400 6 wb_clk_i
port 38 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 42500 42500
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 5203538
string GDS_FILE /run/media/tholin/fbc90f8f-67e9-406d-9872-54f02ad6a2d8/AS2650/openlane/timers/runs/23_11_18_01_08/results/signoff/timers.magic.gds
string GDS_START 439076
<< end >>

