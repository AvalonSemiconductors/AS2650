VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sid_top
  CLASS BLOCK ;
  FOREIGN sid_top ;
  ORIGIN 0.000 0.000 ;
  SIZE 750.000 BY 750.000 ;
  PIN DAC_clk
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 13.440 746.000 14.000 750.000 ;
    END
  END DAC_clk
  PIN DAC_dat_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 64.960 746.000 65.520 750.000 ;
    END
  END DAC_dat_1
  PIN DAC_dat_2
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 90.720 746.000 91.280 750.000 ;
    END
  END DAC_dat_2
  PIN DAC_le
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 39.200 746.000 39.760 750.000 ;
    END
  END DAC_le
  PIN addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 116.480 746.000 117.040 750.000 ;
    END
  END addr[0]
  PIN addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 142.240 746.000 142.800 750.000 ;
    END
  END addr[1]
  PIN addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 168.000 746.000 168.560 750.000 ;
    END
  END addr[2]
  PIN addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 193.760 746.000 194.320 750.000 ;
    END
  END addr[3]
  PIN addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 219.520 746.000 220.080 750.000 ;
    END
  END addr[4]
  PIN bus_cyc
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 657.440 746.000 658.000 750.000 ;
    END
  END bus_cyc
  PIN bus_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 245.280 746.000 245.840 750.000 ;
    END
  END bus_in[0]
  PIN bus_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 271.040 746.000 271.600 750.000 ;
    END
  END bus_in[1]
  PIN bus_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 296.800 746.000 297.360 750.000 ;
    END
  END bus_in[2]
  PIN bus_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 322.560 746.000 323.120 750.000 ;
    END
  END bus_in[3]
  PIN bus_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 348.320 746.000 348.880 750.000 ;
    END
  END bus_in[4]
  PIN bus_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 374.080 746.000 374.640 750.000 ;
    END
  END bus_in[5]
  PIN bus_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 399.840 746.000 400.400 750.000 ;
    END
  END bus_in[6]
  PIN bus_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 425.600 746.000 426.160 750.000 ;
    END
  END bus_in[7]
  PIN bus_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 451.360 746.000 451.920 750.000 ;
    END
  END bus_out[0]
  PIN bus_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 477.120 746.000 477.680 750.000 ;
    END
  END bus_out[1]
  PIN bus_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 502.880 746.000 503.440 750.000 ;
    END
  END bus_out[2]
  PIN bus_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 528.640 746.000 529.200 750.000 ;
    END
  END bus_out[3]
  PIN bus_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 554.400 746.000 554.960 750.000 ;
    END
  END bus_out[4]
  PIN bus_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 580.160 746.000 580.720 750.000 ;
    END
  END bus_out[5]
  PIN bus_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 605.920 746.000 606.480 750.000 ;
    END
  END bus_out[6]
  PIN bus_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 631.680 746.000 632.240 750.000 ;
    END
  END bus_out[7]
  PIN bus_we
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 683.200 746.000 683.760 750.000 ;
    END
  END bus_we
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.738000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 708.960 746.000 709.520 750.000 ;
    END
  END clk
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 734.720 746.000 735.280 750.000 ;
    END
  END rst
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 22.240 15.380 23.840 733.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 15.380 177.440 733.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 329.440 15.380 331.040 733.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 483.040 15.380 484.640 733.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 636.640 15.380 638.240 733.340 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 99.040 15.380 100.640 733.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 252.640 15.380 254.240 733.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 406.240 15.380 407.840 733.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 559.840 15.380 561.440 733.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 713.440 15.380 715.040 733.340 ;
    END
  END vss
  OBS
      LAYER Nwell ;
        RECT 6.290 730.880 743.550 733.470 ;
      LAYER Pwell ;
        RECT 6.290 727.360 743.550 730.880 ;
      LAYER Nwell ;
        RECT 6.290 727.235 63.880 727.360 ;
        RECT 6.290 723.165 743.550 727.235 ;
        RECT 6.290 723.040 37.905 723.165 ;
      LAYER Pwell ;
        RECT 6.290 719.520 743.550 723.040 ;
      LAYER Nwell ;
        RECT 6.290 719.395 19.425 719.520 ;
        RECT 6.290 715.325 743.550 719.395 ;
        RECT 6.290 715.200 12.705 715.325 ;
      LAYER Pwell ;
        RECT 6.290 711.680 743.550 715.200 ;
      LAYER Nwell ;
        RECT 6.290 711.555 62.200 711.680 ;
        RECT 6.290 707.485 743.550 711.555 ;
        RECT 6.290 707.360 333.800 707.485 ;
      LAYER Pwell ;
        RECT 6.290 703.840 743.550 707.360 ;
      LAYER Nwell ;
        RECT 6.290 703.715 91.105 703.840 ;
        RECT 6.290 699.645 743.550 703.715 ;
        RECT 6.290 699.520 12.705 699.645 ;
      LAYER Pwell ;
        RECT 6.290 696.000 743.550 699.520 ;
      LAYER Nwell ;
        RECT 6.290 695.875 142.065 696.000 ;
        RECT 6.290 691.805 743.550 695.875 ;
        RECT 6.290 691.680 12.705 691.805 ;
      LAYER Pwell ;
        RECT 6.290 688.160 743.550 691.680 ;
      LAYER Nwell ;
        RECT 6.290 688.035 105.320 688.160 ;
        RECT 6.290 683.965 743.550 688.035 ;
        RECT 6.290 683.840 149.905 683.965 ;
      LAYER Pwell ;
        RECT 6.290 680.320 743.550 683.840 ;
      LAYER Nwell ;
        RECT 6.290 680.195 12.705 680.320 ;
        RECT 6.290 676.125 743.550 680.195 ;
        RECT 6.290 676.000 39.350 676.125 ;
      LAYER Pwell ;
        RECT 6.290 672.480 743.550 676.000 ;
      LAYER Nwell ;
        RECT 6.290 672.355 22.830 672.480 ;
        RECT 6.290 668.285 743.550 672.355 ;
        RECT 6.290 668.160 81.030 668.285 ;
      LAYER Pwell ;
        RECT 6.290 664.640 743.550 668.160 ;
      LAYER Nwell ;
        RECT 6.290 664.515 180.145 664.640 ;
        RECT 6.290 660.445 743.550 664.515 ;
        RECT 6.290 660.320 14.990 660.445 ;
      LAYER Pwell ;
        RECT 6.290 656.800 743.550 660.320 ;
      LAYER Nwell ;
        RECT 6.290 656.675 36.915 656.800 ;
        RECT 6.290 652.605 743.550 656.675 ;
        RECT 6.290 652.480 38.230 652.605 ;
      LAYER Pwell ;
        RECT 6.290 648.960 743.550 652.480 ;
      LAYER Nwell ;
        RECT 6.290 648.835 25.910 648.960 ;
        RECT 6.290 644.765 743.550 648.835 ;
        RECT 6.290 644.640 51.670 644.765 ;
      LAYER Pwell ;
        RECT 6.290 641.120 743.550 644.640 ;
      LAYER Nwell ;
        RECT 6.290 640.995 140.040 641.120 ;
        RECT 6.290 636.925 743.550 640.995 ;
        RECT 6.290 636.800 12.705 636.925 ;
      LAYER Pwell ;
        RECT 6.290 633.280 743.550 636.800 ;
      LAYER Nwell ;
        RECT 6.290 633.155 185.960 633.280 ;
        RECT 6.290 629.085 743.550 633.155 ;
        RECT 6.290 628.960 32.305 629.085 ;
      LAYER Pwell ;
        RECT 6.290 625.440 743.550 628.960 ;
      LAYER Nwell ;
        RECT 6.290 625.315 12.705 625.440 ;
        RECT 6.290 621.245 743.550 625.315 ;
        RECT 6.290 621.120 51.000 621.245 ;
      LAYER Pwell ;
        RECT 6.290 617.600 743.550 621.120 ;
      LAYER Nwell ;
        RECT 6.290 617.475 144.520 617.600 ;
        RECT 6.290 613.405 743.550 617.475 ;
        RECT 6.290 613.280 83.590 613.405 ;
      LAYER Pwell ;
        RECT 6.290 609.760 743.550 613.280 ;
      LAYER Nwell ;
        RECT 6.290 609.635 18.385 609.760 ;
        RECT 6.290 605.565 743.550 609.635 ;
        RECT 6.290 605.440 21.210 605.565 ;
      LAYER Pwell ;
        RECT 6.290 601.920 743.550 605.440 ;
      LAYER Nwell ;
        RECT 6.290 601.795 56.430 601.920 ;
        RECT 6.290 597.725 743.550 601.795 ;
        RECT 6.290 597.600 74.955 597.725 ;
      LAYER Pwell ;
        RECT 6.290 594.080 743.550 597.600 ;
      LAYER Nwell ;
        RECT 6.290 593.955 38.085 594.080 ;
        RECT 6.290 589.885 743.550 593.955 ;
        RECT 6.290 589.760 81.175 589.885 ;
      LAYER Pwell ;
        RECT 6.290 586.240 743.550 589.760 ;
      LAYER Nwell ;
        RECT 6.290 586.115 9.995 586.240 ;
        RECT 6.290 582.045 743.550 586.115 ;
        RECT 6.290 581.920 55.310 582.045 ;
      LAYER Pwell ;
        RECT 6.290 578.400 743.550 581.920 ;
      LAYER Nwell ;
        RECT 6.290 578.275 136.680 578.400 ;
        RECT 6.290 574.205 743.550 578.275 ;
        RECT 6.290 574.080 39.630 574.205 ;
      LAYER Pwell ;
        RECT 6.290 570.560 743.550 574.080 ;
      LAYER Nwell ;
        RECT 6.290 570.435 27.030 570.560 ;
        RECT 6.290 566.365 743.550 570.435 ;
        RECT 6.290 566.240 80.230 566.365 ;
      LAYER Pwell ;
        RECT 6.290 562.720 743.550 566.240 ;
      LAYER Nwell ;
        RECT 6.290 562.595 57.830 562.720 ;
        RECT 6.290 558.525 743.550 562.595 ;
        RECT 6.290 558.400 204.440 558.525 ;
      LAYER Pwell ;
        RECT 6.290 554.880 743.550 558.400 ;
      LAYER Nwell ;
        RECT 6.290 554.755 130.865 554.880 ;
        RECT 6.290 550.685 743.550 554.755 ;
        RECT 6.290 550.560 110.705 550.685 ;
      LAYER Pwell ;
        RECT 6.290 547.040 743.550 550.560 ;
      LAYER Nwell ;
        RECT 6.290 546.915 224.945 547.040 ;
        RECT 6.290 542.845 743.550 546.915 ;
        RECT 6.290 542.720 48.310 542.845 ;
      LAYER Pwell ;
        RECT 6.290 539.200 743.550 542.720 ;
      LAYER Nwell ;
        RECT 6.290 539.075 222.705 539.200 ;
        RECT 6.290 535.005 743.550 539.075 ;
        RECT 6.290 534.880 21.990 535.005 ;
      LAYER Pwell ;
        RECT 6.290 531.360 743.550 534.880 ;
      LAYER Nwell ;
        RECT 6.290 531.235 150.465 531.360 ;
        RECT 6.290 527.165 743.550 531.235 ;
        RECT 6.290 527.040 203.880 527.165 ;
      LAYER Pwell ;
        RECT 6.290 523.520 743.550 527.040 ;
      LAYER Nwell ;
        RECT 6.290 523.395 12.705 523.520 ;
        RECT 6.290 519.325 743.550 523.395 ;
        RECT 6.290 519.200 71.505 519.325 ;
      LAYER Pwell ;
        RECT 6.290 515.680 743.550 519.200 ;
      LAYER Nwell ;
        RECT 6.290 515.555 18.305 515.680 ;
        RECT 6.290 511.485 743.550 515.555 ;
        RECT 6.290 511.360 12.705 511.485 ;
      LAYER Pwell ;
        RECT 6.290 507.840 743.550 511.360 ;
      LAYER Nwell ;
        RECT 6.290 507.715 92.785 507.840 ;
        RECT 6.290 503.645 743.550 507.715 ;
        RECT 6.290 503.520 165.025 503.645 ;
      LAYER Pwell ;
        RECT 6.290 500.000 743.550 503.520 ;
      LAYER Nwell ;
        RECT 6.290 499.875 34.545 500.000 ;
        RECT 6.290 495.805 743.550 499.875 ;
        RECT 6.290 495.680 86.950 495.805 ;
      LAYER Pwell ;
        RECT 6.290 492.160 743.550 495.680 ;
      LAYER Nwell ;
        RECT 6.290 492.035 21.105 492.160 ;
        RECT 6.290 487.965 743.550 492.035 ;
        RECT 6.290 487.840 12.705 487.965 ;
      LAYER Pwell ;
        RECT 6.290 484.320 743.550 487.840 ;
      LAYER Nwell ;
        RECT 6.290 484.195 142.625 484.320 ;
        RECT 6.290 480.125 743.550 484.195 ;
        RECT 6.290 480.000 159.425 480.125 ;
      LAYER Pwell ;
        RECT 6.290 476.480 743.550 480.000 ;
      LAYER Nwell ;
        RECT 6.290 476.355 90.740 476.480 ;
        RECT 6.290 472.285 743.550 476.355 ;
        RECT 6.290 472.160 12.705 472.285 ;
      LAYER Pwell ;
        RECT 6.290 468.640 743.550 472.160 ;
      LAYER Nwell ;
        RECT 6.290 468.515 52.230 468.640 ;
        RECT 6.290 464.445 743.550 468.515 ;
        RECT 6.290 464.320 40.900 464.445 ;
      LAYER Pwell ;
        RECT 6.290 460.800 743.550 464.320 ;
      LAYER Nwell ;
        RECT 6.290 460.675 39.115 460.800 ;
        RECT 6.290 456.605 743.550 460.675 ;
        RECT 6.290 456.480 42.475 456.605 ;
      LAYER Pwell ;
        RECT 6.290 452.960 743.550 456.480 ;
      LAYER Nwell ;
        RECT 6.290 452.835 170.625 452.960 ;
        RECT 6.290 448.765 743.550 452.835 ;
        RECT 6.290 448.640 12.705 448.765 ;
      LAYER Pwell ;
        RECT 6.290 445.120 743.550 448.640 ;
      LAYER Nwell ;
        RECT 6.290 444.995 61.515 445.120 ;
        RECT 6.290 440.925 743.550 444.995 ;
        RECT 6.290 440.800 110.705 440.925 ;
      LAYER Pwell ;
        RECT 6.290 437.280 743.550 440.800 ;
      LAYER Nwell ;
        RECT 6.290 437.155 111.590 437.280 ;
        RECT 6.290 433.085 743.550 437.155 ;
        RECT 6.290 432.960 83.480 433.085 ;
      LAYER Pwell ;
        RECT 6.290 429.440 743.550 432.960 ;
      LAYER Nwell ;
        RECT 6.290 429.315 12.705 429.440 ;
        RECT 6.290 425.245 743.550 429.315 ;
        RECT 6.290 425.120 153.825 425.245 ;
      LAYER Pwell ;
        RECT 6.290 421.600 743.550 425.120 ;
      LAYER Nwell ;
        RECT 6.290 421.475 56.945 421.600 ;
        RECT 6.290 417.405 743.550 421.475 ;
        RECT 6.290 417.280 187.505 417.405 ;
      LAYER Pwell ;
        RECT 6.290 413.760 743.550 417.280 ;
      LAYER Nwell ;
        RECT 6.290 413.635 287.105 413.760 ;
        RECT 6.290 409.565 743.550 413.635 ;
        RECT 6.290 409.440 41.890 409.565 ;
      LAYER Pwell ;
        RECT 6.290 405.920 743.550 409.440 ;
      LAYER Nwell ;
        RECT 6.290 405.795 12.705 405.920 ;
        RECT 6.290 401.725 743.550 405.795 ;
        RECT 6.290 401.600 154.385 401.725 ;
      LAYER Pwell ;
        RECT 6.290 398.080 743.550 401.600 ;
      LAYER Nwell ;
        RECT 6.290 397.955 12.705 398.080 ;
        RECT 6.290 393.885 743.550 397.955 ;
        RECT 6.290 393.760 29.010 393.885 ;
      LAYER Pwell ;
        RECT 6.290 390.240 743.550 393.760 ;
      LAYER Nwell ;
        RECT 6.290 390.115 38.555 390.240 ;
        RECT 6.290 386.045 743.550 390.115 ;
        RECT 6.290 385.920 36.830 386.045 ;
      LAYER Pwell ;
        RECT 6.290 382.400 743.550 385.920 ;
      LAYER Nwell ;
        RECT 6.290 382.275 209.265 382.400 ;
        RECT 6.290 378.205 743.550 382.275 ;
        RECT 6.290 378.080 112.385 378.205 ;
      LAYER Pwell ;
        RECT 6.290 374.560 743.550 378.080 ;
      LAYER Nwell ;
        RECT 6.290 374.435 12.705 374.560 ;
        RECT 6.290 370.365 743.550 374.435 ;
        RECT 6.290 370.240 76.940 370.365 ;
      LAYER Pwell ;
        RECT 6.290 366.720 743.550 370.240 ;
      LAYER Nwell ;
        RECT 6.290 366.595 52.860 366.720 ;
        RECT 6.290 362.525 743.550 366.595 ;
        RECT 6.290 362.400 13.265 362.525 ;
      LAYER Pwell ;
        RECT 6.290 358.880 743.550 362.400 ;
      LAYER Nwell ;
        RECT 6.290 358.755 110.360 358.880 ;
        RECT 6.290 354.685 743.550 358.755 ;
        RECT 6.290 354.560 209.825 354.685 ;
      LAYER Pwell ;
        RECT 6.290 351.040 743.550 354.560 ;
      LAYER Nwell ;
        RECT 6.290 350.915 130.070 351.040 ;
        RECT 6.290 346.845 743.550 350.915 ;
        RECT 6.290 346.720 335.305 346.845 ;
      LAYER Pwell ;
        RECT 6.290 343.200 743.550 346.720 ;
      LAYER Nwell ;
        RECT 6.290 343.075 12.705 343.200 ;
        RECT 6.290 339.005 743.550 343.075 ;
        RECT 6.290 338.880 13.265 339.005 ;
      LAYER Pwell ;
        RECT 6.290 335.360 743.550 338.880 ;
      LAYER Nwell ;
        RECT 6.290 335.235 98.385 335.360 ;
        RECT 6.290 331.165 743.550 335.235 ;
        RECT 6.290 331.040 160.760 331.165 ;
      LAYER Pwell ;
        RECT 6.290 327.520 743.550 331.040 ;
      LAYER Nwell ;
        RECT 6.290 327.395 218.875 327.520 ;
        RECT 6.290 323.325 743.550 327.395 ;
        RECT 6.290 323.200 88.520 323.325 ;
      LAYER Pwell ;
        RECT 6.290 319.680 743.550 323.200 ;
      LAYER Nwell ;
        RECT 6.290 319.555 16.065 319.680 ;
        RECT 6.290 315.485 743.550 319.555 ;
        RECT 6.290 315.360 12.705 315.485 ;
      LAYER Pwell ;
        RECT 6.290 311.840 743.550 315.360 ;
      LAYER Nwell ;
        RECT 6.290 311.715 32.305 311.840 ;
        RECT 6.290 307.645 743.550 311.715 ;
        RECT 6.290 307.520 91.990 307.645 ;
      LAYER Pwell ;
        RECT 6.290 304.000 743.550 307.520 ;
      LAYER Nwell ;
        RECT 6.290 303.875 24.465 304.000 ;
        RECT 6.290 299.805 743.550 303.875 ;
        RECT 6.290 299.680 45.745 299.805 ;
      LAYER Pwell ;
        RECT 6.290 296.160 743.550 299.680 ;
      LAYER Nwell ;
        RECT 6.290 296.035 62.545 296.160 ;
        RECT 6.290 291.965 743.550 296.035 ;
        RECT 6.290 291.840 44.105 291.965 ;
      LAYER Pwell ;
        RECT 6.290 288.320 743.550 291.840 ;
      LAYER Nwell ;
        RECT 6.290 288.195 16.950 288.320 ;
        RECT 6.290 284.125 743.550 288.195 ;
        RECT 6.290 284.000 59.020 284.125 ;
      LAYER Pwell ;
        RECT 6.290 280.480 743.550 284.000 ;
      LAYER Nwell ;
        RECT 6.290 280.355 51.670 280.480 ;
        RECT 6.290 276.285 743.550 280.355 ;
        RECT 6.290 276.160 149.905 276.285 ;
      LAYER Pwell ;
        RECT 6.290 272.640 743.550 276.160 ;
      LAYER Nwell ;
        RECT 6.290 272.515 36.375 272.640 ;
        RECT 6.290 268.445 743.550 272.515 ;
        RECT 6.290 268.320 159.260 268.445 ;
      LAYER Pwell ;
        RECT 6.290 264.800 743.550 268.320 ;
      LAYER Nwell ;
        RECT 6.290 264.675 256.455 264.800 ;
        RECT 6.290 260.605 743.550 264.675 ;
        RECT 6.290 260.480 201.190 260.605 ;
      LAYER Pwell ;
        RECT 6.290 256.960 743.550 260.480 ;
      LAYER Nwell ;
        RECT 6.290 256.835 29.550 256.960 ;
        RECT 6.290 252.765 743.550 256.835 ;
        RECT 6.290 252.640 9.950 252.765 ;
      LAYER Pwell ;
        RECT 6.290 249.120 743.550 252.640 ;
      LAYER Nwell ;
        RECT 6.290 248.995 166.210 249.120 ;
        RECT 6.290 244.925 743.550 248.995 ;
        RECT 6.290 244.800 158.865 244.925 ;
      LAYER Pwell ;
        RECT 6.290 241.280 743.550 244.800 ;
      LAYER Nwell ;
        RECT 6.290 241.155 37.950 241.280 ;
        RECT 6.290 237.085 743.550 241.155 ;
        RECT 6.290 236.960 154.650 237.085 ;
      LAYER Pwell ;
        RECT 6.290 233.440 743.550 236.960 ;
      LAYER Nwell ;
        RECT 6.290 233.315 51.670 233.440 ;
        RECT 6.290 229.245 743.550 233.315 ;
        RECT 6.290 229.120 210.430 229.245 ;
      LAYER Pwell ;
        RECT 6.290 225.600 743.550 229.120 ;
      LAYER Nwell ;
        RECT 6.290 225.475 48.590 225.600 ;
        RECT 6.290 221.405 743.550 225.475 ;
        RECT 6.290 221.280 62.870 221.405 ;
      LAYER Pwell ;
        RECT 6.290 217.760 743.550 221.280 ;
      LAYER Nwell ;
        RECT 6.290 217.635 413.990 217.760 ;
        RECT 6.290 213.565 743.550 217.635 ;
        RECT 6.290 213.440 227.275 213.565 ;
      LAYER Pwell ;
        RECT 6.290 209.920 743.550 213.440 ;
      LAYER Nwell ;
        RECT 6.290 209.795 186.910 209.920 ;
        RECT 6.290 205.725 743.550 209.795 ;
        RECT 6.290 205.600 86.390 205.725 ;
      LAYER Pwell ;
        RECT 6.290 202.080 743.550 205.600 ;
      LAYER Nwell ;
        RECT 6.290 201.955 138.750 202.080 ;
        RECT 6.290 197.885 743.550 201.955 ;
        RECT 6.290 197.760 41.870 197.885 ;
      LAYER Pwell ;
        RECT 6.290 194.240 743.550 197.760 ;
      LAYER Nwell ;
        RECT 6.290 194.115 118.590 194.240 ;
        RECT 6.290 190.045 743.550 194.115 ;
        RECT 6.290 189.920 177.390 190.045 ;
      LAYER Pwell ;
        RECT 6.290 186.400 743.550 189.920 ;
      LAYER Nwell ;
        RECT 6.290 186.275 11.675 186.400 ;
        RECT 6.290 182.205 743.550 186.275 ;
        RECT 6.290 182.080 28.990 182.205 ;
      LAYER Pwell ;
        RECT 6.290 178.560 743.550 182.080 ;
      LAYER Nwell ;
        RECT 6.290 178.435 89.505 178.560 ;
        RECT 6.290 174.365 743.550 178.435 ;
        RECT 6.290 174.240 68.190 174.365 ;
      LAYER Pwell ;
        RECT 6.290 170.720 743.550 174.240 ;
      LAYER Nwell ;
        RECT 6.290 170.595 22.830 170.720 ;
        RECT 6.290 166.525 743.550 170.595 ;
        RECT 6.290 166.400 245.990 166.525 ;
      LAYER Pwell ;
        RECT 6.290 162.880 743.550 166.400 ;
      LAYER Nwell ;
        RECT 6.290 162.755 259.435 162.880 ;
        RECT 6.290 158.685 743.550 162.755 ;
        RECT 6.290 158.560 12.750 158.685 ;
      LAYER Pwell ;
        RECT 6.290 155.040 743.550 158.560 ;
      LAYER Nwell ;
        RECT 6.290 154.915 9.435 155.040 ;
        RECT 6.290 150.845 743.550 154.915 ;
        RECT 6.290 150.720 47.470 150.845 ;
      LAYER Pwell ;
        RECT 6.290 147.200 743.550 150.720 ;
      LAYER Nwell ;
        RECT 6.290 147.075 67.630 147.200 ;
        RECT 6.290 143.005 743.550 147.075 ;
        RECT 6.290 142.880 51.390 143.005 ;
      LAYER Pwell ;
        RECT 6.290 139.360 743.550 142.880 ;
      LAYER Nwell ;
        RECT 6.290 139.235 260.550 139.360 ;
        RECT 6.290 135.165 743.550 139.235 ;
        RECT 6.290 135.040 59.790 135.165 ;
      LAYER Pwell ;
        RECT 6.290 131.520 743.550 135.040 ;
      LAYER Nwell ;
        RECT 6.290 131.395 79.390 131.520 ;
        RECT 6.290 127.325 743.550 131.395 ;
        RECT 6.290 127.200 18.350 127.325 ;
      LAYER Pwell ;
        RECT 6.290 123.680 743.550 127.200 ;
      LAYER Nwell ;
        RECT 6.290 123.555 35.990 123.680 ;
        RECT 6.290 119.485 743.550 123.555 ;
        RECT 6.290 119.360 31.790 119.485 ;
      LAYER Pwell ;
        RECT 6.290 115.840 743.550 119.360 ;
      LAYER Nwell ;
        RECT 6.290 115.715 14.990 115.840 ;
        RECT 6.290 111.645 743.550 115.715 ;
        RECT 6.290 111.520 40.540 111.645 ;
      LAYER Pwell ;
        RECT 6.290 108.000 743.550 111.520 ;
      LAYER Nwell ;
        RECT 6.290 107.875 16.460 108.000 ;
        RECT 6.290 103.805 743.550 107.875 ;
        RECT 6.290 103.680 33.750 103.805 ;
      LAYER Pwell ;
        RECT 6.290 100.160 743.550 103.680 ;
      LAYER Nwell ;
        RECT 6.290 100.035 14.990 100.160 ;
        RECT 6.290 95.965 743.550 100.035 ;
        RECT 6.290 95.840 107.950 95.965 ;
      LAYER Pwell ;
        RECT 6.290 92.320 743.550 95.840 ;
      LAYER Nwell ;
        RECT 6.290 92.195 32.350 92.320 ;
        RECT 6.290 88.125 743.550 92.195 ;
        RECT 6.290 88.000 23.670 88.125 ;
      LAYER Pwell ;
        RECT 6.290 84.480 743.550 88.000 ;
      LAYER Nwell ;
        RECT 6.290 84.355 52.300 84.480 ;
        RECT 6.290 80.285 743.550 84.355 ;
        RECT 6.290 80.160 50.865 80.285 ;
      LAYER Pwell ;
        RECT 6.290 76.640 743.550 80.160 ;
      LAYER Nwell ;
        RECT 6.290 76.515 43.270 76.640 ;
        RECT 6.290 72.445 743.550 76.515 ;
        RECT 6.290 72.320 51.435 72.445 ;
      LAYER Pwell ;
        RECT 6.290 68.800 743.550 72.320 ;
      LAYER Nwell ;
        RECT 6.290 68.675 35.990 68.800 ;
        RECT 6.290 64.605 743.550 68.675 ;
        RECT 6.290 64.480 157.275 64.605 ;
      LAYER Pwell ;
        RECT 6.290 60.960 743.550 64.480 ;
      LAYER Nwell ;
        RECT 6.290 60.835 54.680 60.960 ;
        RECT 6.290 56.765 743.550 60.835 ;
        RECT 6.290 56.640 68.190 56.765 ;
      LAYER Pwell ;
        RECT 6.290 53.120 743.550 56.640 ;
      LAYER Nwell ;
        RECT 6.290 52.995 43.270 53.120 ;
        RECT 6.290 48.925 743.550 52.995 ;
        RECT 6.290 48.800 74.955 48.925 ;
      LAYER Pwell ;
        RECT 6.290 45.280 743.550 48.800 ;
      LAYER Nwell ;
        RECT 6.290 45.155 51.670 45.280 ;
        RECT 6.290 41.085 743.550 45.155 ;
        RECT 6.290 40.960 110.785 41.085 ;
      LAYER Pwell ;
        RECT 6.290 37.440 743.550 40.960 ;
      LAYER Nwell ;
        RECT 6.290 37.315 62.590 37.440 ;
        RECT 6.290 33.245 743.550 37.315 ;
        RECT 6.290 33.120 123.420 33.245 ;
      LAYER Pwell ;
        RECT 6.290 29.600 743.550 33.120 ;
      LAYER Nwell ;
        RECT 6.290 29.475 76.310 29.600 ;
        RECT 6.290 25.405 743.550 29.475 ;
        RECT 6.290 25.280 116.630 25.405 ;
      LAYER Pwell ;
        RECT 6.290 21.760 743.550 25.280 ;
      LAYER Nwell ;
        RECT 6.290 21.635 193.690 21.760 ;
        RECT 6.290 17.440 743.550 21.635 ;
      LAYER Pwell ;
        RECT 6.290 15.250 743.550 17.440 ;
      LAYER Metal1 ;
        RECT 6.720 15.380 743.120 734.570 ;
      LAYER Metal2 ;
        RECT 6.860 745.700 13.140 746.000 ;
        RECT 14.300 745.700 38.900 746.000 ;
        RECT 40.060 745.700 64.660 746.000 ;
        RECT 65.820 745.700 90.420 746.000 ;
        RECT 91.580 745.700 116.180 746.000 ;
        RECT 117.340 745.700 141.940 746.000 ;
        RECT 143.100 745.700 167.700 746.000 ;
        RECT 168.860 745.700 193.460 746.000 ;
        RECT 194.620 745.700 219.220 746.000 ;
        RECT 220.380 745.700 244.980 746.000 ;
        RECT 246.140 745.700 270.740 746.000 ;
        RECT 271.900 745.700 296.500 746.000 ;
        RECT 297.660 745.700 322.260 746.000 ;
        RECT 323.420 745.700 348.020 746.000 ;
        RECT 349.180 745.700 373.780 746.000 ;
        RECT 374.940 745.700 399.540 746.000 ;
        RECT 400.700 745.700 425.300 746.000 ;
        RECT 426.460 745.700 451.060 746.000 ;
        RECT 452.220 745.700 476.820 746.000 ;
        RECT 477.980 745.700 502.580 746.000 ;
        RECT 503.740 745.700 528.340 746.000 ;
        RECT 529.500 745.700 554.100 746.000 ;
        RECT 555.260 745.700 579.860 746.000 ;
        RECT 581.020 745.700 605.620 746.000 ;
        RECT 606.780 745.700 631.380 746.000 ;
        RECT 632.540 745.700 657.140 746.000 ;
        RECT 658.300 745.700 682.900 746.000 ;
        RECT 684.060 745.700 708.660 746.000 ;
        RECT 709.820 745.700 734.420 746.000 ;
        RECT 735.580 745.700 741.300 746.000 ;
        RECT 6.860 7.370 741.300 745.700 ;
      LAYER Metal3 ;
        RECT 6.810 7.420 741.350 733.180 ;
      LAYER Metal4 ;
        RECT 21.420 15.080 21.940 731.270 ;
        RECT 24.140 15.080 98.740 731.270 ;
        RECT 100.940 15.080 175.540 731.270 ;
        RECT 177.740 15.080 252.340 731.270 ;
        RECT 254.540 15.080 329.140 731.270 ;
        RECT 331.340 15.080 405.940 731.270 ;
        RECT 408.140 15.080 482.740 731.270 ;
        RECT 484.940 15.080 559.540 731.270 ;
        RECT 561.740 15.080 636.340 731.270 ;
        RECT 638.540 15.080 709.940 731.270 ;
        RECT 21.420 7.930 709.940 15.080 ;
  END
END sid_top
END LIBRARY

