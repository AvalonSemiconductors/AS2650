* NGSPICE file created from wrapped_as2650.ext - technology: gf180mcuC

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__antenna abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__antenna I VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_1 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_1 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_64 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_64 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_1 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_2 I0 I1 S Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_1 D CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_4 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__tiel abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__tiel ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_2 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__tieh abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__tieh Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_2 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_1 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_4 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_2 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_1 A1 A2 A3 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_1 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_1 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_2 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_1 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_2 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_1 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_1 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_1 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi222_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_1 A1 A2 B1 B2 C1 C2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor3_2 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_2 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_2 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_2 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_2 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_1 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux4_2 I0 I1 I2 I3 S0 S1 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_2 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_4 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_1 A1 A2 A3 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_4 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_4 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_4 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_2 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_1 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyc_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyc_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi222_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_4 A1 A2 B1 B2 C1 C2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_2 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyb_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyb_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_4 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_2 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_1 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_2 D CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_2 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_2 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_4 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_2 A1 A2 A3 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_4 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_4 A1 A2 A3 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_4 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux4_1 I0 I1 I2 I3 S0 S1 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_2 A1 A2 A3 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai33_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai33_1 A1 A2 A3 B1 B2 B3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi222_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_2 A1 A2 B1 B2 C1 C2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux4_4 I0 I1 I2 I3 S0 S1 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai222_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai222_2 A1 A2 B1 B2 C1 C2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_2 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai222_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai222_1 A1 A2 B1 B2 C1 C2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_2 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_2 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_2 A1 A2 A3 Z VDD VSS
.ends

.subckt wrapped_as2650 io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14]
+ io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22]
+ io_in[23] io_in[24] io_in[25] io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30]
+ io_in[31] io_in[32] io_in[33] io_in[34] io_in[35] io_in[36] io_in[37] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_in[8] io_in[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12]
+ io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1]
+ io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27]
+ io_oeb[28] io_oeb[29] io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34]
+ io_oeb[35] io_oeb[36] io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7]
+ io_oeb[8] io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14]
+ io_out[15] io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21]
+ io_out[22] io_out[23] io_out[24] io_out[25] io_out[26] io_out[27] io_out[28] io_out[29]
+ io_out[2] io_out[30] io_out[31] io_out[32] io_out[33] io_out[34] io_out[35] io_out[36]
+ io_out[37] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9]
+ la_data_out[0] la_data_out[10] la_data_out[11] la_data_out[12] la_data_out[13] la_data_out[14]
+ la_data_out[15] la_data_out[16] la_data_out[17] la_data_out[18] la_data_out[19]
+ la_data_out[1] la_data_out[20] la_data_out[21] la_data_out[22] la_data_out[23] la_data_out[24]
+ la_data_out[25] la_data_out[26] la_data_out[27] la_data_out[28] la_data_out[29]
+ la_data_out[2] la_data_out[30] la_data_out[31] la_data_out[32] la_data_out[33] la_data_out[34]
+ la_data_out[35] la_data_out[36] la_data_out[37] la_data_out[38] la_data_out[39]
+ la_data_out[3] la_data_out[40] la_data_out[41] la_data_out[42] la_data_out[43] la_data_out[44]
+ la_data_out[45] la_data_out[46] la_data_out[47] la_data_out[48] la_data_out[49]
+ la_data_out[4] la_data_out[50] la_data_out[51] la_data_out[52] la_data_out[53] la_data_out[54]
+ la_data_out[55] la_data_out[56] la_data_out[57] la_data_out[58] la_data_out[59]
+ la_data_out[5] la_data_out[60] la_data_out[61] la_data_out[62] la_data_out[63] la_data_out[6]
+ la_data_out[7] la_data_out[8] la_data_out[9] vdd vss wb_clk_i
XFILLER_132_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07383__I _01817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05903_ _05756_ _05757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06883_ _01251_ _01303_ _01323_ _01324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09671_ _03787_ _03788_ _03833_ _03834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07534__A1 _01854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05834_ as2650.ins_reg\[1\] _05688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08622_ net94 _02776_ _02894_ _02895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_27_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08553_ _01610_ _02826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_36_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09287__A1 as2650.stack\[2\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_165_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07504_ as2650.stack\[7\]\[13\] _01933_ _01934_ as2650.stack\[6\]\[13\] _01935_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_08484_ _01143_ _02733_ _02757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__07837__A2 _02197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05848__A1 _05700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10841__A1 _04167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07435_ _01791_ _01869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_167_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09039__A1 _01884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10249__I _03165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07366_ _01801_ _01802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_182_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09105_ _05731_ _01358_ _03328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06317_ _00766_ _00767_ _00768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_104_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07297_ _01732_ _01733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_178_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09036_ _03265_ as2650.r123_2\[0\]\[1\] _03259_ _03266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06248_ _00679_ _00574_ _00704_ _00705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_164_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06812__A3 _01253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_1861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_191_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_163_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06179_ _00637_ _00638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_172_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06025__A1 net72 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07222__B1 _01658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08565__A3 _05793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09762__A2 _03920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07773__A1 _02122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11812__CLK clknet_leaf_111_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09938_ _00717_ _04094_ _02890_ _04095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_104_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07293__I net48 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_189_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09869_ _01465_ _01457_ _04027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_100_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11900_ _00269_ clknet_leaf_73_wb_clk_i as2650.stack\[6\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output37_I net37 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11962__CLK clknet_leaf_20_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11831_ _00214_ clknet_leaf_27_wb_clk_i as2650.r123_2\[1\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_165_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08338__B _02640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_104_wb_clk_i_I clknet_4_3_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10587__C _04643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11762_ _00145_ clknet_leaf_82_wb_clk_i as2650.stack\[5\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10713_ _01737_ _04822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10832__A1 _03639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11693_ _00076_ clknet_leaf_119_wb_clk_i as2650.stack\[11\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09948__I _00957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10644_ _03921_ _03964_ _04754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_167_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_155_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10575_ _02789_ _04685_ _04686_ _04687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_13_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09450__A1 as2650.stack\[5\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08253__A2 _00834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06372__I _00817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07461__B1 _01863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07461__C2 as2650.stack\[1\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08005__A2 _02357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06016__A1 _05678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07764__A1 _02177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11127_ _01811_ _05225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_122_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09505__A2 _03669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11058_ _01942_ _05157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_67_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06319__A2 _00646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07516__A1 as2650.stack\[9\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11312__A2 _05268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10009_ _02893_ _04165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_49_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_168_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10778__B _03641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09269__A1 _03475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11076__A1 as2650.stack\[10\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_181_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11076__B2 as2650.stack\[8\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10823__A1 _00627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_177_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08492__A2 _02726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07220_ _01628_ _01656_ _01657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_20_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_34_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11379__A2 _05457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07151_ _01166_ _01567_ _01579_ _01588_ _01589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_125_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08244__A2 _00483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09441__A1 as2650.stack\[5\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_146_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10587__B1 _04680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06102_ as2650.cycle\[5\] _00561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_157_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06282__I _00735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07082_ _05775_ _01362_ _01521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_195_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_173_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06033_ _00463_ _00492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__11835__CLK clknet_leaf_32_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_173_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06007__A1 _05728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10960__C _00786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11000__A1 _01091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08547__A3 _01430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09744__A2 _03901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07755__A1 _02078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11551__A2 _05140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10532__I _04404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07984_ _02347_ _02352_ _02353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_87_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11985__CLK clknet_leaf_77_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05861__S0 _05685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09723_ _03836_ _03837_ _03884_ _03885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08002__I _02073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06935_ _01373_ _01361_ _01374_ _01375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_132_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07507__A1 as2650.stack\[5\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11303__A2 _05302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07507__B2 as2650.stack\[4\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09654_ _00805_ _00816_ _03817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06866_ _01027_ _01307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_27_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10511__B1 _01794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xwrapped_as2650_104 io_oeb[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_08605_ _01406_ _01490_ _02878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_27_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05817_ _05670_ _05671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xwrapped_as2650_115 io_out[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_06797_ _01187_ _01191_ _01176_ _01239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_09585_ _02865_ _03749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_27_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_126 la_data_out[35] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_55_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_137 la_data_out[56] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xwrapped_as2650_148 io_oeb[34] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XTAP_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11067__A1 as2650.stack\[2\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08536_ _02808_ _02809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xwrapped_as2650_159 la_data_out[46] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XANTENNA__11067__B2 as2650.stack\[0\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10200__C _04349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10814__A1 _04913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08467_ _00964_ _02740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09680__A1 _03796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08483__A2 _02755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06494__A1 _00459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07418_ as2650.r123\[0\]\[2\] _01852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08398_ _02236_ _02686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_91_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07349_ as2650.stack\[11\]\[8\] _01740_ _01784_ _01785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08235__A2 _02530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10578__B1 _04681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07288__I _01723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10360_ _00881_ _00979_ _04482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__06192__I _05728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07994__A1 _01984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09019_ _03249_ _03250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_151_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10291_ _02332_ _02847_ _04427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_3_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12030_ _00399_ clknet_leaf_51_wb_clk_i as2650.r123\[3\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_137_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06549__A2 _00544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07746__A1 as2650.stack\[11\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11542__A2 _02153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_43_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_115_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08171__A1 _02321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_185_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06721__A2 _01127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11814_ _00197_ clknet_leaf_108_wb_clk_i as2650.stack\[1\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_163_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11745_ _00128_ clknet_4_8_0_wb_clk_i as2650.stack\[7\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_42_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07277__A3 _00963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08582__I _02854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11676_ _00059_ clknet_leaf_128_wb_clk_i as2650.stack\[13\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_35_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_146_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11858__CLK clknet_leaf_32_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10627_ as2650.stack\[13\]\[3\] _01751_ _02795_ as2650.stack\[12\]\[3\] _04738_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_139_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11230__A1 _05129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10558_ _01271_ _05754_ _04670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_128_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_155_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07985__B2 _00853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10489_ _04585_ _04589_ _04594_ _04601_ _04602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_48_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06830__I _01271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06720_ _01133_ _01153_ _01162_ _01055_ _01163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__08162__A1 _02133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06651_ _01082_ _01085_ _01089_ _01094_ _01095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_64_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_111_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06582_ _00930_ _00612_ _01026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09370_ _03561_ _03562_ _03563_ _03564_ _00263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06277__I _00730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08321_ as2650.stack\[4\]\[8\] _02627_ _02629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09662__A1 _03824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08465__A2 _00542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09588__I _03751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08252_ _00605_ _00798_ _00873_ _02555_ _02561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XANTENNA__10272__A2 _04309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07203_ _05723_ _01109_ _01640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_177_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08183_ _02186_ _02485_ _02486_ _02506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__10527__I _03915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08217__A2 _02491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09414__A1 _03571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_192_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06228__A1 _00524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07134_ _01568_ _00666_ _01571_ _01572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_88_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11221__A1 _00757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09965__A2 _04120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_134_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07065_ _01352_ _01369_ _01386_ _01503_ _01504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_145_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10690__C _04798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07836__I _02046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09029__S _03259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06016_ _05678_ _00446_ _00452_ _00474_ _00475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XANTENNA__12013__CLK clknet_leaf_106_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09717__A2 _03878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07991__A4 _02023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07728__A1 _02143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06400__A1 _00831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07967_ _00837_ _00464_ _02335_ _02336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_114_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09706_ _03836_ _03867_ _00679_ _03868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06918_ _01358_ _01359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_28_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07898_ _02051_ _02270_ _02283_ _02287_ _00068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__07571__I _01991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09637_ _03798_ _03799_ _03800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06849_ _00957_ _01291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10211__B _04103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07900__A1 _02167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09568_ net93 _03732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_110_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08519_ _02789_ _02790_ _02791_ _02792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_130_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09499_ _00929_ _03665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_51_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06467__A1 _00694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10865__C _02809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11530_ _05557_ _05577_ _05578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10263__A2 _02606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11461_ _02901_ _02844_ _05521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__09405__A1 _03561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10015__A2 _02940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10412_ _02553_ _03598_ _04526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__11212__A1 as2650.stack\[14\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11392_ as2650.stack\[9\]\[13\] _05464_ _05470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__11212__B2 as2650.stack\[12\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10343_ _04467_ _00333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_124_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10274_ _00978_ _00822_ _04412_ _04413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_140_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07719__A1 _02133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11515__A2 _02770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12013_ _00382_ clknet_leaf_106_wb_clk_i as2650.stack\[9\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_120_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08577__I _02849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08144__A1 _02321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09892__A1 _03957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09892__B2 _02105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06097__I _00555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05902__B1 _05754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11680__CLK clknet_leaf_131_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_159_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06458__A1 as2650.cycle\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_175_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10254__A2 _04392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11728_ _00111_ clknet_leaf_115_wb_clk_i as2650.stack\[0\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_9_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10347__I _04469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11659_ _00042_ clknet_leaf_126_wb_clk_i as2650.stack\[11\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_106_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_174_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11203__A1 as2650.stack\[6\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11203__B2 as2650.stack\[4\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07958__A1 _02327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07656__I _02080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11506__A2 _04463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08870_ _01142_ _03082_ _03115_ _03116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_111_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10714__B1 _01793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07821_ _02222_ _02227_ _02228_ _02210_ _00050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_111_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10190__A1 _00863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06933__A2 _01198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10810__I _04595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07752_ as2650.stack\[11\]\[3\] _02149_ _02169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_96_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05904__I as2650.r0\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08135__A1 _02153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07391__I _01825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06703_ _00433_ _00435_ _01146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07683_ _02105_ _02106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_20_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09422_ _03603_ _00276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06634_ _01031_ _01074_ _01078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_53_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09353_ _02284_ _02658_ _03551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06565_ as2650.idx_ctrl\[0\] _01009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09635__A1 _01041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08438__A2 _02707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_4_5_0_wb_clk_i_I clknet_3_2_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08304_ _02612_ _02613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_21_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06496_ _05714_ _00940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09284_ _03020_ _03494_ _03497_ _03498_ _00243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_20_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08235_ as2650.stack\[5\]\[14\] _02530_ _02545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_176_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06464__A4 _00581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_193_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09938__A2 _04094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08166_ _02487_ _02495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_194_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07949__A1 _02321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_194_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07117_ _01376_ _01548_ _01554_ _01512_ _01555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_134_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08097_ _02418_ _02442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08171__B _02494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07048_ as2650.holding_reg\[5\] _01486_ _01483_ _01487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_122_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_102_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07177__A2 _01614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08374__A1 as2650.stack\[2\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_134_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08999_ _02097_ _03222_ _03234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_125_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08126__A1 as2650.stack\[0\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09323__B1 _03525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_117_wb_clk_i clknet_4_2_0_wb_clk_i clknet_leaf_117_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_44_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_84_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10961_ _00784_ _00681_ _05062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_16_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09874__A1 _04025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06688__A1 _00541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10484__A2 as2650.ins_reg\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10892_ _01884_ _04995_ _04979_ _03667_ _00882_ _04996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_58_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08429__A2 _02491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11433__A1 _01137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09021__I _03249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11513_ _01306_ _00859_ _05192_ _02608_ _05562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_184_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06860__A1 _01008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11444_ _05508_ _05509_ _00392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08860__I _03103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11375_ as2650.stack\[9\]\[8\] _05456_ _05458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_180_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08081__B _02424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06380__I _00477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10326_ _04454_ _00783_ _00786_ _04340_ _04455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_112_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10257_ _00976_ _04400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09905__B _04062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07168__A2 _01605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08365__A1 as2650.stack\[3\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10188_ _00563_ _02547_ _04338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_61_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10172__A1 _02561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08117__A1 _02405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10786__B _04887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06350_ _00798_ _00799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_148_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11424__A1 _03568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_187_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_104_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06281_ _00734_ _00735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_30_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09866__I _00534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08020_ _02128_ _02381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_163_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10805__I _00711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06603__A1 _00428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09971_ _04124_ _04126_ _04127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08922_ _01436_ _03165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_131_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout86_I net59 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08853_ _00606_ _00745_ _01024_ _03100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_97_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10163__A1 _00808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10540__I _04651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07804_ _02213_ _02214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_61_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08784_ _03033_ _03022_ _03034_ _03036_ _00205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_85_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05996_ _00447_ _00455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__08108__A1 _02399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07735_ _02154_ _02137_ _02034_ _02155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XTAP_2908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09856__A1 _04000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_187_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07666_ _02089_ _02090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_168_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07331__A2 _01747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09405_ _03561_ _03589_ _03590_ _03591_ _00271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06617_ as2650.holding_reg\[0\] _01061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_13_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07597_ _02024_ _02025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07882__A3 _02147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06465__I _00466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09336_ _03044_ _03533_ _03536_ _03537_ _00256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06548_ _00743_ _00992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_139_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09267_ _03477_ _03479_ _03483_ _03484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_166_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06479_ _00922_ _00923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_166_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08680__I _02932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08218_ _02533_ _02534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11919__CLK clknet_leaf_96_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09198_ _03416_ _03417_ _03418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_105_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08149_ as2650.stack\[8\]\[12\] _02477_ _02482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_88_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08595__A1 _02834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07398__A2 _01832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11160_ _01747_ _05257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07229__C _01486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10111_ _04256_ _04099_ _03727_ _04264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_161_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11091_ _05124_ _05189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_5501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_136_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10042_ _02205_ _04069_ _04196_ _04163_ _04197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA_output67_I net67 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10154__A1 _03699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_5545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_102_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_102_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06373__A3 _00818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09847__A1 _03977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11993_ _00362_ clknet_leaf_19_wb_clk_i as2650.r0\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_57_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10457__A2 _00687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10944_ _04255_ _04270_ _04988_ _05046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_28_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10875_ _02211_ _04974_ _04979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_16_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08076__B _02424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_38_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xclkbuf_leaf_85_wb_clk_i clknet_4_2_0_wb_clk_i clknet_leaf_85_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XPHY_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07086__A1 _05732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12029__D _00398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_185_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_160_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08804__B _03021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06833__A1 _01274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_51_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09619__C _03782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11427_ _03571_ _05487_ _05494_ _05495_ _00389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_137_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11358_ as2650.r123_2\[3\]\[1\] _05448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_152_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10309_ _04426_ _04441_ _04442_ _00324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_11289_ _05238_ _04081_ _05382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_141_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08338__A1 _02521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10145__A1 _02225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10145__B2 _00452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05850_ _05700_ _05704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_55_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09838__A1 net35 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_99_wb_clk_i_I clknet_4_9_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07520_ _01766_ _01949_ _01950_ _01951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_47_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08765__I _01983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08510__A1 as2650.stack\[7\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07313__A2 _01729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08510__B2 as2650.stack\[6\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07451_ _01263_ _01803_ _01885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_23_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06402_ _00842_ _00847_ _00848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_34_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05875__A2 _05728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07382_ _01755_ _01817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09121_ _03303_ _03335_ _03343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_148_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06333_ _00782_ _00783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08813__A2 _03055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09596__I _00722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06824__A1 _01265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06264_ _00718_ _00719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09052_ _01927_ _03279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_124_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09529__C _03692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08003_ _02368_ _02365_ _02369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06195_ _00653_ _00654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09954_ _02808_ _04008_ _04111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08329__A1 _02513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08905_ _01309_ _03149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09885_ _04041_ _04042_ _04043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__10136__A1 _04270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10136__B2 net92 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11333__B1 _03679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10270__I _03991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07001__A1 _01431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08836_ _01043_ _03082_ _03083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09541__A3 _02572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06355__A3 _00770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08767_ _03021_ _03022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09829__A1 _02612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05979_ _00424_ _05785_ _00422_ _00438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_122_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07718_ _01988_ _02138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10439__A2 _04552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08698_ _02709_ _02969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08501__A1 _00853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07649_ _02036_ _02074_ _02063_ _02075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_14_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_40_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_148_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06195__I _00653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10660_ _04766_ _04768_ _04769_ _04588_ _04770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_16_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11741__CLK clknet_leaf_116_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09319_ _02284_ _02639_ _03525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_90_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_161_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10591_ _02081_ _04646_ _04702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__07607__A3 _02034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06815__A1 _01008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_194_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_107_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11891__CLK clknet_leaf_94_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11212_ as2650.stack\[14\]\[3\] _05268_ _05269_ as2650.stack\[12\]\[3\] _05215_ _05308_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_147_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput20 net20 io_oeb[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput31 net31 io_out[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput42 net42 io_out[32] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_11143_ _00775_ _01249_ _05237_ _05239_ _05240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_134_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput53 net94 la_data_out[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput64 net88 la_data_out[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_163_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput75 net75 la_data_out[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_163_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07791__A2 _02202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_132_wb_clk_i clknet_4_0_0_wb_clk_i clknet_leaf_132_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_163_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_133_wb_clk_i_I clknet_4_1_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10127__A1 _03759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11074_ as2650.stack\[9\]\[0\] _05171_ _05172_ as2650.stack\[11\]\[0\] _05173_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_5331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10127__B2 _03772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11324__B1 _05414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10025_ _03794_ _04177_ _04179_ _03769_ _04180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_49_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_5364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05929__I0 as2650.r123\[1\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09532__A3 _00870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10678__A2 _04748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06346__A3 _00684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08740__A1 _02384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08740__B2 _03002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_149_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_188_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11627__A1 _02616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08585__I _01436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11976_ _00345_ clknet_leaf_75_wb_clk_i net56 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10927_ _00794_ _04293_ _05029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_17_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10858_ _04226_ _04946_ _04963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10850__A2 _04192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_157_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10789_ _02902_ _04889_ _04895_ _04819_ _04896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XPHY_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_118_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06806__A1 _01082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10602__A2 _04711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06806__B2 _01077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_184_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08559__A1 _02813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_172_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10366__A1 net43 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07231__A1 _01666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_101_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06951_ _01390_ _01167_ _01391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11186__I _00680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05902_ _05752_ _05726_ _05754_ _05718_ _05755_ _05706_ _05756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_132_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09670_ _03814_ _03831_ _03832_ _03833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06882_ _01305_ _01315_ _01322_ _01154_ _01250_ _01323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__09523__A3 _03686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08731__A1 _02415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08621_ _02893_ _02894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05833_ net54 _05687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_94_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08552_ _01598_ _02590_ _02822_ _02824_ _02825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__11618__A1 _05413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08495__I _02583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11764__CLK clknet_leaf_94_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05912__I _05765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07503_ _01824_ _01934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_36_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08483_ _02754_ _02755_ _02756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07434_ _01864_ _01867_ _01846_ _01868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_195_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_51_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07365_ _01105_ _01710_ _01801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_149_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08444__B _02718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09104_ as2650.r0\[6\] _01217_ _03327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_149_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06316_ _05704_ _00590_ _00767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_52_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07296_ _01731_ _01732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_148_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09035_ _03129_ _03245_ _03248_ _03264_ _03265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__10265__I _04404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06247_ _00702_ _00703_ _00704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_117_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06178_ as2650.addr_buff\[7\] _00637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10357__A1 _04326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_1884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07222__A1 as2650.r123\[1\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_85_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09275__B _03489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08565__A4 _02837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07574__I _01819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08970__A1 _02345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07773__A2 _02172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09937_ _04092_ _04093_ _04094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_131_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11306__B1 _05257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06981__B1 _01420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09868_ _01609_ _01618_ _04026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11029__C _03781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07525__A2 _01953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08722__A1 as2650.stack\[15\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08819_ _00987_ _00995_ _03054_ _03066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XTAP_3214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09722__C _03883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09799_ _03879_ _03959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_189_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11830_ _00213_ clknet_leaf_33_wb_clk_i as2650.r123_2\[1\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11609__A1 _01290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06918__I _01358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11609__B2 _05647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05822__I _05675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_27_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11761_ _00144_ clknet_leaf_82_wb_clk_i as2650.stack\[5\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11085__A2 _05183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_158_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10712_ _04237_ _04817_ _04820_ _04821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_1878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10832__A2 _04934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11692_ _00075_ clknet_leaf_119_wb_clk_i as2650.stack\[11\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_41_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10643_ _04654_ _04749_ _04751_ _04752_ _04753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_195_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07749__I _02073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_158_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10574_ as2650.stack\[2\]\[2\] _04681_ _02914_ as2650.stack\[0\]\[2\] _04686_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__10596__A1 _00446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09450__A2 _03615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08073__C _02424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10175__I _02608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07461__A1 as2650.stack\[3\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_182_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11637__CLK clknet_leaf_36_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06016__A2 _00446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08961__A1 _01589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07764__A2 _02178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11126_ as2650.stack\[9\]\[1\] _02142_ _05223_ as2650.stack\[11\]\[1\] _05224_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_68_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11057_ _01940_ _05156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_5161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11787__CLK clknet_leaf_85_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07516__A2 _01942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08713__A1 _02449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10008_ _02195_ _04069_ _04162_ _04163_ _04164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XTAP_5194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10520__A1 _04626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07433__B _01866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09269__A2 _03484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_51_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11076__A2 _01959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11959_ _00328_ clknet_4_5_0_wb_clk_i as2650.holding_reg\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_177_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10823__A2 _05721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_189_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08492__A3 _02727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07150_ _01327_ _01584_ _01587_ _01588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_125_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_173_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09441__A2 _03615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_185_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06101_ _00458_ _00557_ _00559_ _00560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_07081_ _01514_ _01519_ _01520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_161_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06032_ _05691_ _00491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_138_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06007__A2 _00465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11000__A2 _02723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08547__A4 _01265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07394__I _01828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08952__A1 _05801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11551__A3 _02768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07983_ _02351_ _02352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_59_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09722_ _02071_ _03725_ _03882_ _03883_ _03884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_06934_ _05760_ _01109_ _01374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05861__S1 _05714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10969__B _02331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08704__A1 _02276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07507__A2 _01936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09901__B1 _00817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09653_ _02608_ _03816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06865_ _01265_ _01306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09542__C _03705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10511__A1 as2650.stack\[6\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10511__B2 as2650.stack\[4\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05908__I3 as2650.r123_2\[0\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08604_ _01420_ _01412_ _01480_ _01488_ _02877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08180__A2 _02488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05816_ _05669_ _05670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_27_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xwrapped_as2650_105 io_oeb[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_09584_ _03740_ _00683_ _03742_ _03732_ _03747_ _03748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_3_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xwrapped_as2650_116 io_out[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_06796_ _01237_ _01238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_127 la_data_out[37] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08535_ _02807_ _02808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_24_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xwrapped_as2650_138 la_data_out[58] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xwrapped_as2650_149 io_oeb[35] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XANTENNA__11067__A2 _01940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10814__A2 _04077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08466_ _00867_ _02583_ _02738_ _00849_ _02739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_195_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07417_ _01807_ _01720_ _01851_ _00023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_11_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06494__A2 _00937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08397_ _02684_ _02681_ _02682_ _02685_ _00169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_11_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07569__I _01996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_177_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07348_ _01765_ _01784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_6_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10578__A1 as2650.stack\[11\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10578__B2 as2650.stack\[10\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07279_ _00947_ _00953_ _01305_ _01007_ _01715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_164_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09018_ _01725_ _03101_ _03249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_139_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07994__A2 _02357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10290_ _04425_ _04426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_2_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05817__I _05670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08943__A1 _01474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07746__A2 _02163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10750__A1 _01697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10502__A1 _00689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08171__A2 _02489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06182__A1 _00540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_160_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11813_ _00196_ clknet_leaf_111_wb_clk_i as2650.stack\[1\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11744_ _00127_ clknet_leaf_114_wb_clk_i as2650.stack\[8\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09671__A2 _03788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07277__A4 _01712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_169_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11675_ _00058_ clknet_leaf_128_wb_clk_i as2650.stack\[13\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_169_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07479__I _01717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10626_ as2650.stack\[15\]\[3\] _02782_ _01780_ as2650.stack\[14\]\[3\] _04737_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_127_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07434__A1 _01864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10557_ net10 _05754_ _04669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_122_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11230__A2 _02223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05928__S _05753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10488_ _04596_ _04582_ _04600_ _04432_ _04601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_139_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11518__B1 _05565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09187__A1 _03145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10633__I _04529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10741__A1 _01465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_4_12_0_wb_clk_i clknet_3_6_0_wb_clk_i clknet_4_12_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_11109_ _04460_ _03679_ _05204_ _03782_ _05206_ _05207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_42_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09643__B _01002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08162__A2 _02491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06558__I _00961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06650_ _01093_ _01094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_77_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06581_ _00745_ _01024_ _00942_ _01025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_18_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08320_ _02627_ _02628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_162_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08251_ _00785_ _02549_ _02559_ _02560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_33_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07389__I _01823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07202_ _01637_ _01638_ _01639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_20_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06293__I _00744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08182_ _02196_ _02505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08217__A3 _02471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09414__A2 _03589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07133_ _01569_ _00962_ _01570_ _00666_ _01571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__06228__A2 _00685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11221__A2 _05294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10971__C _04554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07064_ _01214_ _01353_ _01366_ _01385_ _01503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_118_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11952__CLK clknet_4_5_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06015_ _00473_ _00474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07338__B net73 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08925__A1 _01599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07728__A2 _02146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_192_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_99_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08013__I _02109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07966_ _00503_ _01087_ _02335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09705_ _03866_ _03867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06917_ as2650.r123\[0\]\[3\] as2650.r123_2\[0\]\[3\] _05709_ _01358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11288__A2 _05381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07897_ _02284_ _02285_ _02286_ _02287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09350__A1 _02045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09636_ _03796_ _01118_ _01158_ _03799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
X_06848_ _01103_ _01290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06468__I _00774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09567_ _03729_ _03730_ _03731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_71_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06779_ _01215_ _01220_ _01221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_130_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08518_ as2650.stack\[2\]\[6\] _01745_ _01756_ as2650.stack\[0\]\[6\] _02791_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08683__I _01697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09498_ _03636_ _03660_ _03664_ _00697_ _00291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_93_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10799__A1 _04237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11323__B _00914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07664__A1 _02078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08449_ _05670_ _02722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_157_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07664__B2 _02088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07299__I _01734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11460_ _02616_ _05520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__11042__C _05140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09405__A2 _03589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07416__A1 _01808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10411_ _00637_ _02013_ _04341_ _04525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_139_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11212__A2 _05268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11391_ _02680_ _05467_ _05468_ _05469_ _00379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_10_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07967__A2 _00464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10342_ _04399_ _04463_ _04458_ _00827_ _04467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_109_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_152_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09169__A1 _03366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10971__A1 _00783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10971__B2 _04364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10273_ _03706_ _04408_ _04410_ _04411_ _04412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_3_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09019__I _03249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12012_ _00381_ clknet_4_2_0_wb_clk_i as2650.stack\[9\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_45_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_155_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10723__A1 _02789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_leaf_39_wb_clk_i clknet_4_6_0_wb_clk_i clknet_leaf_39_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_132_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08858__I _03104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07762__I _02109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08079__B _02424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08144__A2 _02468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09341__A1 _02129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06378__I _00823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06155__A1 _00492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_185_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09892__A2 net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05902__A1 _05752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05902__B2 _05718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11825__CLK clknet_leaf_100_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06458__A2 _00561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11727_ _00110_ clknet_leaf_88_wb_clk_i as2650.stack\[0\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_159_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11658_ _00041_ clknet_leaf_124_wb_clk_i as2650.stack\[11\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11975__CLK clknet_leaf_75_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10609_ _04669_ _04673_ _04719_ _04720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__07407__A1 _01765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08604__B1 _01480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11203__A2 _05296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09801__C1 _00818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11589_ _02746_ _00951_ _05633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_176_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07958__A2 _02279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05969__A1 _05773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10962__A1 _01155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_123_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10714__A1 as2650.stack\[7\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10714__B2 as2650.stack\[4\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07820_ as2650.stack\[14\]\[12\] _02208_ _02228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09373__B _03543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06394__A1 _00503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10190__A2 _02722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07751_ _02067_ _02141_ _02166_ _02168_ _00040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_187_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06702_ _01144_ _01145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_38_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08135__A2 _01989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09332__A1 _02456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07682_ net61 _02105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_37_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09421_ as2650.ivec\[1\] _03261_ _03601_ _03603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06633_ _00884_ _00515_ _01077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_129_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09599__I _03762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09352_ _02049_ _03550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_178_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06564_ _00960_ _01008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_52_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09635__A2 _01018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08303_ _02611_ _02612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_94_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07646__A1 _01263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11442__A2 _03406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09283_ _03000_ _02673_ _02682_ _03498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__10538__I _04649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06495_ _00646_ _00938_ _00939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08234_ _02525_ _02541_ _02542_ _02544_ _00147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_165_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_165_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_140_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09399__A1 as2650.stack\[6\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08165_ _02314_ _02489_ _02490_ _02494_ _00128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_88_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07116_ _05751_ _01360_ _01510_ _01357_ _01554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_147_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_140_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08096_ as2650.stack\[0\]\[0\] _02440_ _02441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_133_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10953__A1 _05026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07068__B _01361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07047_ _01228_ _01486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_134_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10705__A1 _00978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09571__A1 _03732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09283__B _02682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06385__A1 _05696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08998_ _02493_ _03233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_75_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07949_ _02321_ _02315_ _02322_ _02317_ _00084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_75_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08126__A2 _02445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09323__A1 _03028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10960_ _04811_ _05057_ _05060_ _00786_ _05061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_112_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06688__A2 _00812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09619_ _03775_ _03778_ _03780_ _03782_ _03783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_16_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10891_ _04622_ _04995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_188_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05830__I _05683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07637__A1 as2650.stack\[13\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11512_ _00826_ _00846_ _05561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_157_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11443_ _01295_ _05502_ _05504_ as2650.r123\[2\]\[2\] _05509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06860__A2 _01009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09458__B _03621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_153_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11374_ _05456_ _05457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_193_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10944__A1 _04255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10325_ _04376_ _04454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_49_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06612__A2 _01019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10256_ _02861_ _04399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_152_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08365__A2 _02655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08588__I _02826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10187_ net91 _04337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_121_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10172__A2 _02563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08117__A2 _02454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11121__A1 _05216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07876__A1 _02237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_72_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11424__A2 _05487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10632__B1 _04741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06280_ as2650.cycle\[8\] _00734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06300__A1 _00707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_175_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11188__A1 _03761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07667__I _02090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08053__A1 _02405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_171_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09970_ _03849_ _04125_ _04126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07800__A1 _02189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08921_ _03110_ _03162_ _03164_ _00214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_130_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08852_ _00921_ _03067_ _03099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_44_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06367__A1 _00720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_131_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10163__A2 _00608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07803_ _01219_ _02191_ _02192_ _02212_ _02213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_08783_ as2650.stack\[8\]\[2\] _03035_ _03031_ _03036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05995_ _00453_ _05692_ _00454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08108__A2 _02436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09305__A1 as2650.stack\[2\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07734_ _02153_ _02154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_72_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06119__A1 _00480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07665_ _00940_ _02089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09404_ as2650.stack\[6\]\[4\] _03585_ _03582_ _03591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06616_ net50 net78 _01060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07596_ _01999_ _02001_ _02003_ _02023_ _02024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_146_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09335_ _02989_ _02634_ _03518_ _03537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_142_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06547_ _00990_ _00991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09266_ _03480_ _03482_ _03483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_142_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06478_ _00491_ _00898_ _00922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08292__B2 _00753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08217_ _01985_ _02491_ _02471_ _02533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_193_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06842__A2 _01157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09197_ _03397_ _03398_ _03417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__11179__A1 _05265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08148_ _02473_ _02481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08044__A1 _02399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10926__A1 _05026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08595__A2 _00769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08079_ _02321_ _02420_ _02424_ _02428_ _00108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_84_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_162_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09792__I net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10110_ _03867_ _04262_ _04263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11090_ _03974_ _05188_ _00359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_81_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_clkbuf_leaf_123_wb_clk_i_I clknet_4_2_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09544__A1 _05703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10041_ _04185_ _04195_ _04196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_5524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_102_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06358__A1 _00805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05825__I as2650.ins_reg\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11351__A1 _05221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_5579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_188_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_4845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12026__CLK clknet_leaf_39_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11103__A1 _04275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11992_ _00361_ clknet_4_5_0_wb_clk_i as2650.r0\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_28_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_56_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09847__A2 _02890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10887__B _04363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_186_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10943_ _04242_ _04988_ _04395_ _05045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_72_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06656__I _01022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10874_ _04223_ _03733_ _04977_ _04978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_44_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06530__A1 net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09032__I _03249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_157_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07086__A2 _01109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_184_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_61_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10090__A1 _04242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_145_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06391__I _05685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11426_ as2650.stack\[9\]\[7\] _05476_ _05472_ _05495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_86_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10917__A1 _03755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_54_wb_clk_i clknet_4_13_0_wb_clk_i clknet_leaf_54_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_125_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09783__A1 _02853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11357_ _05447_ _00367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_152_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09916__B _03887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11590__A1 _00662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05939__A4 _05769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10308_ as2650.holding_reg\[3\] _04423_ _04442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_158_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11288_ _05281_ _05381_ _00364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_3_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09535__A1 _00852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10239_ _04385_ _04387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10145__A2 _04111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11342__A1 _05430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07010__A2 _01449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09550__A4 _00956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07950__I _02219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07849__A1 as2650.stack\[13\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08510__A2 _02782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07450_ _01861_ _01868_ _01882_ _01883_ _01884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_63_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_179_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06521__A1 _00964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06401_ _00843_ _00846_ _00847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_147_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07381_ _01815_ _01816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_176_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09120_ _03339_ _03342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06332_ _00458_ _00782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08274__A1 _00863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09051_ _03247_ _03278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_148_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10081__A1 _03737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06263_ _00714_ _00718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_163_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07397__I _01810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08002_ _02073_ _02368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_191_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06194_ as2650.ins_reg\[2\] as2650.ins_reg\[3\] _00653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_102_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10908__A1 _04654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_191_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_171_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06588__A1 _01028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11581__A1 _02956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08730__B _02969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09953_ _04098_ _04100_ _04108_ _04109_ _04110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_103_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09526__A1 _03688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08904_ _01234_ _03148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_170_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09884_ _03975_ _03996_ _04042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10136__A2 _04103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11333__A1 _01029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11333__B2 _00810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08835_ _03081_ _03082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_170_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08766_ _02472_ _03021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05978_ _05769_ _00437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_57_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input11_I io_in[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09829__A2 _01474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07717_ _02136_ _02137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08697_ _02905_ _02967_ _02968_ _00186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_26_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08177__B _02501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08501__A2 _02768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06476__I net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07648_ _02073_ _02074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06512__A1 _00645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07579_ _00513_ _00626_ _02007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_15_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10447__I0 _02038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09318_ _03020_ _03519_ _03522_ _03524_ _00251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08265__A1 _05670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10590_ _04700_ _04701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_166_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08624__C _02352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_194_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_166_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09249_ _03419_ _03466_ _03441_ _03442_ _03467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__06815__A2 _01009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08017__A1 as2650.stack\[14\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_194_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11211_ as2650.stack\[13\]\[3\] _05266_ _05172_ as2650.stack\[15\]\[3\] _05307_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_135_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09765__A1 _00689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06579__A1 _01022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput21 net21 io_out[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_162_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11572__A1 _05138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput32 net32 io_out[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_122_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput43 net43 io_out[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_11142_ _05238_ _01286_ _00914_ _05239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_150_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput54 net54 la_data_out[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput65 net87 la_data_out[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__09517__A1 _02726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput76 net76 la_data_out[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_122_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11073_ _01819_ _05172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_5321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10127__A2 _04276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11324__A1 _00775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06160__B _00618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10024_ _04174_ _04178_ _04179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_7_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05929__I1 as2650.r123\[0\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09532__A4 _02555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_5387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08740__A2 _02996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08866__I _03077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_4675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06751__A1 _01166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_101_wb_clk_i clknet_4_3_0_wb_clk_i clknet_leaf_101_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_63_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11627__A2 _04443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11975_ _00344_ clknet_leaf_75_wb_clk_i net55 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08087__B _02431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10926_ _05026_ _05027_ _05028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_166_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10857_ _04157_ _04930_ _04186_ _04962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_108_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09697__I _02889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08256__A1 _02560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10788_ _04651_ _04878_ _04895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_12_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_185_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_160_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_121_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07464__C1 as2650.stack\[10\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08008__A1 _02078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09056__I0 _03282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08106__I _02073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11409_ as2650.stack\[9\]\[2\] _05478_ _05483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_177_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11563__A1 _00471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06950_ _05763_ _01390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_98_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_171_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07519__B1 _01819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input3_I io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05901_ as2650.r123\[1\]\[2\] as2650.r123\[0\]\[2\] as2650.r123_2\[1\]\[2\] as2650.r123_2\[0\]\[2\]
+ _05705_ _05753_ _05755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_132_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06881_ _01317_ _01321_ _01322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_132_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08620_ _00677_ _02893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05832_ _05682_ _05685_ _05686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_95_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08731__A2 _02985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09381__B _03543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11909__CLK clknet_leaf_75_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08551_ _02823_ _02824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__11618__A2 _04638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_184_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07502_ _01836_ _01933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_93_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08482_ _00952_ _00899_ _01986_ _00606_ _02755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06296__I _00485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07433_ as2650.stack\[2\]\[10\] _01865_ _01866_ _01867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_74_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10974__C _04744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07364_ _01760_ _01778_ _01798_ _01799_ _01800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA__08247__A1 _00459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_176_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09103_ _03322_ _03325_ _03326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__10054__A1 _04129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06315_ _05701_ _00766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10054__B2 _04024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07295_ net70 _01730_ _01731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09034_ _03261_ _03262_ _03263_ _03264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06246_ _00544_ _00703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10990__B _03737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06177_ _00635_ _00636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_132_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_85_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08970__A2 _03111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10281__I _02772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09936_ _04049_ _04052_ _04047_ _04093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_120_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11306__A1 as2650.stack\[2\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06981__B2 _01094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11306__B2 as2650.stack\[1\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09867_ _02826_ _04025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_112_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08722__A2 _02978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08818_ _03064_ _03065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06733__A1 as2650.holding_reg\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09798_ _03957_ _03958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_85_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08749_ as2650.stack\[1\]\[3\] _02998_ _03009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_73_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11760_ _00143_ clknet_leaf_81_wb_clk_i as2650.stack\[5\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10293__A1 _01136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10711_ _03642_ _04810_ _04818_ _04819_ _04820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_1857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11691_ _00074_ clknet_leaf_126_wb_clk_i as2650.stack\[10\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_42_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08238__A1 _00992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10642_ _02824_ _04752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_41_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11699__D _00082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10456__I _04225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10573_ as2650.stack\[3\]\[2\] _02908_ _02785_ as2650.stack\[1\]\[2\] _04685_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_195_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10596__A2 _04703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07461__A2 _01862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09738__A1 _03150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11545__A1 _02847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06016__A3 _00452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08410__A1 as2650.stack\[1\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11125_ _01761_ _05223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_123_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_5140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11056_ as2650.stack\[5\]\[0\] _05153_ _05154_ as2650.stack\[7\]\[0\] _05155_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_49_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10007_ _00749_ _04163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08713__A2 _02974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_5184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08477__A1 _00898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11958_ _00327_ clknet_leaf_17_wb_clk_i as2650.holding_reg\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_33_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10284__A1 _00767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10909_ _04391_ _03873_ _05012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_44_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11889_ _00258_ clknet_leaf_102_wb_clk_i as2650.stack\[4\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_149_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08492__A4 _02333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11233__B1 _03679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07437__C1 as2650.stack\[10\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06100_ _00558_ _00559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_34_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07080_ _01020_ _01518_ _01519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_8_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07452__A2 _01884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_173_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09729__A1 _03842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06031_ _00486_ _00489_ _00490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_172_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10339__A2 _00887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11536__A1 _04626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11536__B2 _02621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08401__A1 _02030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08952__A2 _03059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07982_ _02350_ _02351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_138_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11731__CLK clknet_leaf_111_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06933_ _05766_ _01198_ _01373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09721_ _03718_ _03883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09901__A1 _04025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08704__A2 _02974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06864_ _01001_ _00966_ _01128_ _01304_ _01305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__09901__B2 _04041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09652_ _03657_ _03815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_99_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06715__A1 _01120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10511__A2 _01823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05815_ as2650.cycle\[6\] _05669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08603_ _01576_ _01676_ _02876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_27_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09583_ _03732_ _03744_ _03746_ _03747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_82_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06795_ _01233_ _01236_ _01237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_23_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xwrapped_as2650_106 io_oeb[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_97_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xwrapped_as2650_117 io_out[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_83_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08534_ _02806_ _02807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_128 la_data_out[39] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xwrapped_as2650_139 la_data_out[60] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_70_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08468__A1 _05671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08465_ _02582_ _00542_ _02738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_24_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07416_ _01808_ _01722_ _01719_ _01850_ _01851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_195_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_149_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08396_ as2650.stack\[2\]\[13\] _02676_ _02685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_10_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10027__A1 net38 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07347_ as2650.stack\[9\]\[8\] _01762_ _01761_ as2650.stack\[8\]\[8\] as2650.stack\[10\]\[8\]
+ _01782_ _01783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_195_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_176_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10578__A2 _02908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_192_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07278_ _01103_ _01713_ _01052_ _01714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08640__A1 _02907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09017_ _03247_ _03248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06229_ _00562_ _00687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_163_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_1671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_1682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09735__A4 _01285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06954__A1 _01393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10750__A2 _04056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09919_ _04075_ _04076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_output42_I net42 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06706__A1 _01142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05833__I net54 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_189_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11812_ _00195_ clknet_leaf_111_wb_clk_i as2650.stack\[1\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10266__A1 _02778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11743_ _00126_ clknet_leaf_114_wb_clk_i as2650.stack\[8\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_169_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11674_ _00057_ clknet_leaf_132_wb_clk_i as2650.stack\[13\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_109_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11215__B1 _05310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10625_ as2650.stack\[11\]\[3\] _01839_ _02907_ _04736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_122_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09975__I net38 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10556_ _04570_ _04668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_194_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_182_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10487_ _00445_ _04599_ _04600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_6_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11518__A1 _02571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07495__I _01430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06613__B _01056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11518__B2 _02780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09187__A2 _03298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11754__CLK clknet_leaf_81_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07198__A1 as2650.r0\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10741__A2 _05737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11108_ _01146_ _00789_ _05205_ _03138_ _05206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_81_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10789__C _04819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11039_ _00613_ _05138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_64_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08162__A3 _02471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07370__A1 _01721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06580_ _00937_ _01024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_94_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09111__A2 _03333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11480__I _05539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_177_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08250_ _02551_ _02553_ _02556_ _02558_ _02559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__08870__A1 _01142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07201_ _05742_ _01198_ _01638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08181_ _02329_ _02500_ _02501_ _02504_ _00134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_158_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_9_wb_clk_i clknet_4_4_0_wb_clk_i clknet_leaf_9_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07132_ _05748_ _00990_ _01570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__10029__C _00552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08622__A1 net94 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07063_ _01477_ _01501_ _00968_ _01502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_134_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11509__A1 _01992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06014_ _00458_ _00472_ _00473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_47_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08925__A2 _03113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07728__A3 _02147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06936__A1 _01357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07965_ _02333_ _02334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_9_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09704_ _02932_ _03866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06916_ _05780_ _01357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08689__A1 _02960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07896_ _02280_ _02286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_83_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09635_ _01041_ _01018_ _03798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_06847_ _01280_ _01287_ _01288_ _01289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_16_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07361__A1 _01788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06778_ _01020_ _01219_ _01220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09566_ _02037_ _01041_ _03730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_110_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10248__A1 _03150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08517_ as2650.stack\[3\]\[6\] _02782_ _01751_ as2650.stack\[1\]\[6\] _02790_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_130_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09497_ _03662_ _00623_ _03660_ _03663_ _03664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_51_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06484__I _00743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08448_ _02686_ _02717_ _02718_ _02721_ _00184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__07664__A2 _01998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08379_ _02206_ _02672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_71_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_177_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10410_ _00662_ _00704_ _04524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_164_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08613__A1 _01097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11777__CLK clknet_leaf_82_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11390_ as2650.stack\[9\]\[12\] _05464_ _05469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09810__B1 _03916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08632__C _02903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10341_ _00460_ _04457_ _04466_ _00332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__10420__A1 _00799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07967__A3 _02335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05828__I net94 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10272_ _03685_ _04309_ _03689_ _03707_ _04411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XANTENNA__08204__I _02511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12011_ _00380_ clknet_leaf_117_wb_clk_i as2650.stack\[9\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_155_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07719__A3 _02138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06659__I _00955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09341__A2 _02634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06155__A2 _00503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11514__B _05562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11726_ _00109_ clknet_leaf_83_wb_clk_i as2650.stack\[0\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_14_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08852__A1 _00921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_174_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11657_ _00040_ clknet_leaf_124_wb_clk_i as2650.stack\[11\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_156_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10608_ net11 _05767_ _04719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__08604__A1 _01420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11588_ _03642_ _04462_ _02965_ _05632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__09801__C2 _03951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10411__A1 _00637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_183_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10539_ _02350_ _04651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08080__A2 _02427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07439__B _01872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05969__A2 _00427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10962__A2 _05062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07953__I _02226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10714__A2 _04822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06394__A2 _00839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10190__A3 _00627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07174__B _01144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_152_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07750_ _02167_ _02156_ _02164_ _02168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_113_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06701_ _01143_ _01025_ _01144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08135__A3 _02471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09332__A2 _03523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_187_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07681_ _02035_ _02104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_65_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06632_ _01059_ _01075_ _01076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09420_ _03602_ _00275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_64_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06563_ _01001_ _00966_ _01003_ _01006_ _01007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_09351_ _03542_ _03544_ _03547_ _03549_ _00259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_33_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08302_ _01465_ _02611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09282_ as2650.stack\[2\]\[0\] _03496_ _03497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06494_ _00459_ _00937_ _00938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_127_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_166_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08233_ as2650.stack\[5\]\[13\] _02538_ _02544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__10650__A1 _04584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08164_ _02493_ _02494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09399__A2 _03577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_181_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07115_ _05742_ _01108_ _01553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10402__A1 _02551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07349__B _01784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08095_ _02439_ _02440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_173_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06082__A1 _00540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07046_ _01478_ _00667_ _01481_ _01485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_106_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08024__I _01983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_113_wb_clk_i_I clknet_4_2_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_192_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_161_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06909__A1 _01096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_5706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09056__S _03271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10705__A2 _04586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_138_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_134_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09571__A2 _03734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_134_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06385__A2 _00830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08997_ _03037_ _03217_ _03230_ _03232_ _00222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_131_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07582__A1 _00948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06479__I _00922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07948_ as2650.stack\[10\]\[10\] _02319_ _02322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__11318__C _05278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10222__C _03786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07879_ _02269_ _02270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_44_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07334__A1 _01736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09618_ _03781_ _03782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_16_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06688__A3 _01130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10890_ _04948_ _04993_ _04994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09087__A1 _05758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09549_ _00911_ _00574_ _03713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_169_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08834__A1 _01604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07637__A2 _02062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10641__A1 _04596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11511_ _05150_ _05559_ _05560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_133_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_157_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10892__C _00882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11442_ _05496_ _03406_ _05508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_126_wb_clk_i clknet_4_0_0_wb_clk_i clknet_leaf_126_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_166_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11197__A2 _03815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11373_ _05455_ _05456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_158_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10944__A2 _04270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10324_ _04453_ _00328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_3_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_171_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10255_ _04397_ _04388_ _04398_ _00314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_124_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09011__A1 _03050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10186_ net83 _04325_ _04336_ _00307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_120_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10413__B _04308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10172__A3 _02594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06389__I _00834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_187_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_74_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07876__A2 _02263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11942__CLK clknet_leaf_56_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05887__A1 _05735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10639__I _04748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_182_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08825__A1 _00981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10632__A1 _04620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11709_ _00092_ clknet_leaf_0_wb_clk_i as2650.stack\[14\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_147_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06300__A2 _00751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11188__A2 _01303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09250__A1 _01663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08053__A2 _02406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06073__B _00531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10935__A2 _04769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07800__A2 _02207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08920_ _01370_ _03163_ _03130_ as2650.r123_2\[1\]\[3\] _03164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_143_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09002__A1 as2650.stack\[7\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07683__I _02105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08851_ _03069_ _03095_ _03097_ _03098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_150_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09553__A2 _03706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07802_ _02211_ _02212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_69_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06299__I _00750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05994_ _05691_ _00453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08782_ _03025_ _03035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07733_ _02152_ _02153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_84_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06119__A2 _00457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08513__B1 _01756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07867__A2 _02260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07664_ _02078_ _01998_ _02079_ _02088_ _00033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09403_ _03509_ _03579_ _03590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06615_ _01058_ _01059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10871__A1 _04223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07595_ _02022_ _02023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_74_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06546_ _00989_ _00990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_94_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09334_ as2650.stack\[4\]\[5\] _03526_ _03536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_161_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_142_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10993__B _03755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09265_ _03439_ _03443_ _03470_ _03481_ _03482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_06477_ _00851_ _00921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_138_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_166_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07858__I _02255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08216_ as2650.stack\[5\]\[8\] _02530_ _02532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_14_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09196_ _03360_ _03415_ _03416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_194_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11179__A2 _05275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08147_ _02467_ _02480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_159_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08078_ as2650.stack\[0\]\[10\] _02427_ _02428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_49_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_175_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07029_ _01463_ _00933_ _01035_ _01467_ _01468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_121_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__11815__CLK clknet_leaf_111_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07004__B1 _01425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10040_ _02205_ _04111_ _04194_ _03830_ _04195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XTAP_5514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09544__A2 _00458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06358__A2 _00801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11351__A2 _05442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_3_4_0_wb_clk_i_I clknet_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11990__D _00359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11991_ _00360_ clknet_leaf_26_wb_clk_i as2650.r0\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11103__A2 _01127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10942_ _04668_ _05037_ _05039_ _05043_ _05044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_83_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10862__A1 _04879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10873_ _00794_ _04232_ _04977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10862__B2 _04771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06530__A2 _00936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06158__B _00508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09480__A1 _03646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07491__B1 _01900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11425_ _02184_ _05480_ _05494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_153_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06046__A1 _00487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10127__C _03774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11356_ as2650.r123_2\[3\]\[0\] _05447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09783__A2 _03147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10307_ _04438_ _04440_ _04441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_193_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11287_ _03285_ _05189_ _05380_ _05381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_79_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_140_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_94_wb_clk_i clknet_4_10_0_wb_clk_i clknet_leaf_94_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_10238_ _04386_ _00309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_84_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07546__A1 _01975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10143__B _03728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10169_ _00546_ _02599_ _04319_ _04320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_121_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_67_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09424__S _03604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09651__C _03813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09299__A1 _03509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10369__I _04482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_165_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06521__A2 _00926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06400_ _00831_ _00845_ _00846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_37_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07380_ _01814_ _01815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_62_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_76_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_194_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06331_ _00780_ _00781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10605__A1 _04584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08274__A2 _02582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07678__I _02100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09050_ _03277_ _00230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_148_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06285__A1 _00728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06262_ _00551_ _00717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_15_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08001_ _02051_ _02357_ _02363_ _02367_ _00091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_190_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09223__A1 _05724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06193_ _00460_ _00454_ _00652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10908__A2 _05007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06588__A2 _01029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11581__A2 _02609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout91_I net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09952_ _00672_ _04109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_28_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05926__I as2650.r0\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08903_ _01156_ _01298_ _01300_ _01318_ _01320_ _03147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XANTENNA__09526__A2 _03689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08302__I _01465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09883_ net36 _04041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_112_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11333__A2 _02867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08834_ _01604_ _03061_ _03081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_112_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08765_ _01983_ _03020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_85_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05977_ _00428_ _00433_ _00435_ _00436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_100_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11097__A1 _05129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07716_ _02135_ _01993_ _02136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08696_ _02951_ _02776_ _02894_ _02968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_65_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07647_ _02071_ _02041_ _02072_ _02073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_14_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06512__A2 _00558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07578_ _00817_ _02005_ _00956_ _02006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_80_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09317_ _03000_ _03523_ _02640_ _03524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06529_ _00972_ _00973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_178_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09462__A1 _03565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08265__A2 _00735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09248_ _01597_ _03465_ _03466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_127_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08017__A2 _02362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09179_ _03395_ _03399_ _03400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_147_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07076__I0 as2650.r123\[0\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11021__A1 _03646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11210_ _05300_ _05305_ _05222_ _05306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09765__A2 _03903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06579__A2 _00944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput22 net22 io_out[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__11572__A2 _04417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput33 net33 io_out[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_11141_ _00641_ _05238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_134_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput44 net44 io_out[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_150_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput55 net90 la_data_out[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_81_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output72_I net72 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput66 net66 la_data_out[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_1_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09517__A2 _03673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput77 net77 la_data_out[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_11072_ _01812_ _05171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_5300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11324__A2 _01685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10023_ _04156_ _04118_ _04120_ _04178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_118_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_5344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05929__I2 as2650.r123_2\[1\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_5388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11088__A1 _05147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11974_ _00343_ clknet_leaf_49_wb_clk_i net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_56_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10925_ _02217_ _05000_ _05027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_189_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06503__A2 _00946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10856_ _04116_ _04173_ _04930_ _04961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_176_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09453__A1 as2650.stack\[5\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_157_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10787_ _04879_ _04893_ _04894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_13_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07464__B1 _01758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07464__C2 _01747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08008__A2 _02357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09056__I1 as2650.r123_2\[0\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06019__A1 _00476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11012__A1 _00533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_126_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11408_ _03550_ _05473_ _05479_ _05482_ _00383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_114_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11563__A2 _02757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11339_ as2650.stack\[0\]\[7\] _05210_ _05431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08122__I _02118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07519__B2 as2650.stack\[12\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05900_ as2650.r123\[2\]\[2\] as2650.r123_2\[2\]\[2\] _05753_ _05754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_151_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06880_ _01319_ _01300_ _01320_ _01321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_95_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_121_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05831_ _05684_ _05685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_67_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06577__I _01020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08550_ _02607_ _02823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_130_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07501_ _01502_ _01932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_78_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10826__A1 _04668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08481_ _02730_ _02753_ _02754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09692__A1 _03850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07432_ _01734_ _01866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_1_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07363_ _01777_ _01799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08247__A2 _00798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09444__A1 _03542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09444__B2 _03618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09102_ _03320_ _03323_ _03324_ _03325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_148_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06258__A1 _00548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06314_ _00764_ _00765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11251__A1 _05264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07294_ net86 _01729_ _01730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_175_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09033_ _01847_ _03252_ _03263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06245_ _00701_ _00702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_178_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_163_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12016__CLK clknet_leaf_101_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11003__A1 _00864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06176_ _00511_ _00630_ _00633_ _00634_ _00539_ _00635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_102_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_1853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_144_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_1875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11554__A2 _02731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10762__B1 _04845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06430__A1 _00543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09935_ net63 net2 _04092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__08032__I _02250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09866_ _00534_ _04024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10514__B1 _01826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08183__A1 _02186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08817_ _02089_ _00982_ _00967_ _03064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_100_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09797_ net60 _03957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08748_ _02399_ _02996_ _03007_ _03008_ _00197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10817__A1 _04808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08679_ net54 _02951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_41_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09798__I _03957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10710_ _04363_ _04819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10293__A2 _04428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11690_ _00073_ clknet_leaf_0_wb_clk_i as2650.stack\[10\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10641_ _04596_ _04750_ _04751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11342__B _05152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10737__I _04844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08238__A2 _00734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09435__A1 as2650.ivec\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06249__A1 _00700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11242__A1 _05333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07446__B1 _01879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08207__I _02230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08643__C1 as2650.stack\[3\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10572_ _01787_ _04682_ _04683_ _04684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_107_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09738__A2 _03762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_159_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11545__A2 _02770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08410__A2 _02695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09038__I _01263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06421__A1 _00866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11124_ _05151_ _05222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_137_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11055_ _01937_ _05154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_5141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07781__I net88 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10006_ _04135_ _04146_ _04160_ _04161_ _04162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_5174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08098__B _02431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10808__A1 _04875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11957_ _00326_ clknet_leaf_20_wb_clk_i as2650.holding_reg\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_44_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08477__A2 _00598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_181_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10284__A2 _04420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10908_ _04654_ _05007_ _05010_ _04752_ _05011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__11481__A1 _03977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11888_ _00257_ clknet_leaf_102_wb_clk_i as2650.stack\[4\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_127_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09501__I _03666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10839_ _04913_ _04531_ _04944_ _00352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_32_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11233__A1 _03149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07437__B1 _01758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11233__B2 _02860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07437__C2 _01870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07021__I _01390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_179_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06030_ _00488_ _00489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07956__I _02230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_160_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_177_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11536__A2 _05565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08401__A2 _02649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06412__A1 _00824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07981_ _02349_ _02350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_141_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09720_ _03860_ _03869_ _03881_ _00731_ _03882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_101_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06932_ _01352_ _01369_ _01372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_67_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07691__I _02112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08165__A1 _02314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09651_ _03789_ _03792_ _03812_ _03813_ _03814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_132_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09901__A2 _03872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06176__B1 _00634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06863_ _00709_ _00585_ _00642_ _00906_ _01304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_67_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06715__A2 _01156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07912__A1 _02177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08602_ _02874_ _01668_ _02875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_94_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09582_ _03745_ _03746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_55_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06794_ _01234_ _00829_ _01229_ _01235_ _01236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
Xwrapped_as2650_107 io_oeb[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_83_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xwrapped_as2650_118 io_out[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_184_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06100__I _00558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08533_ _00878_ _02806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_110_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_36_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xwrapped_as2650_129 la_data_out[41] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__09665__A1 _02332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08468__A2 _02740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10275__A2 _04412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_3_7_0_wb_clk_i clknet_0_wb_clk_i clknet_3_7_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_24_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08464_ _00950_ _02737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_24_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_168_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07415_ _01728_ _01847_ _01848_ _01849_ _01850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_11_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09417__A1 _03598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08395_ _02230_ _02684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_91_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_195_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11224__A1 _04275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07346_ _01781_ _01782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08027__I _01832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07277_ _00785_ _00974_ _00963_ _01712_ _01713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_104_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09016_ _03102_ _03246_ _03247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__06651__A1 _01082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06228_ _00524_ _00685_ _00686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_164_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10292__I _02349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06159_ _00507_ _00610_ _00617_ _00618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_104_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06954__A2 _00962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09918_ _00626_ _04075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_28_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_clkbuf_leaf_69_wb_clk_i_I clknet_4_9_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09849_ _00800_ _02618_ _04008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_98_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06706__A2 _00934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07903__A1 _02170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output35_I net35 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11811_ _00194_ clknet_leaf_4_wb_clk_i as2650.stack\[15\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_26_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_160_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10895__C _04912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10266__A2 _01024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11742_ _00125_ clknet_leaf_116_wb_clk_i as2650.stack\[8\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11463__A1 _01022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09321__I _02632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11673_ _00056_ clknet_leaf_131_wb_clk_i as2650.stack\[13\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_39_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09408__A1 _03565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11215__A1 as2650.stack\[8\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06890__A1 as2650.holding_reg\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10624_ as2650.stack\[9\]\[3\] _01815_ _01818_ as2650.stack\[8\]\[3\] as2650.stack\[10\]\[3\]
+ _01876_ _04735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_169_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11215__B2 as2650.stack\[11\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10555_ _02902_ _04649_ _04666_ _04667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_154_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07776__I _02187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10486_ _04597_ _04598_ _04599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_4_14_0_wb_clk_i_I clknet_3_7_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_155_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07198__A2 _01378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_151_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11107_ _02745_ _04651_ _05205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_61_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11038_ _05132_ _05133_ _05134_ _05136_ _05137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_37_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09647__A1 net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07200_ _01513_ _01635_ _01636_ _01549_ _01637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_165_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08180_ as2650.stack\[7\]\[14\] _02488_ _02504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_18_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07131_ _05743_ _01569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_140_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08622__A2 _02776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_173_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06590__I _00432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06633__A1 _00884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07062_ _01096_ _01480_ _01494_ _01500_ _01501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_4
XFILLER_122_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06013_ _00459_ _00471_ _00472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_192_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_103_wb_clk_i_I clknet_4_9_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10717__B1 _01825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08386__A1 _02675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_173_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07964_ _02008_ _02333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_87_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08138__A1 _02314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09703_ _03861_ _03864_ _03865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_96_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06915_ _01354_ _01355_ _01356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_114_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_5_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08310__I _02618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09886__A1 _03811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08689__A2 _01700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07895_ _02277_ _02285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09634_ _03796_ _03797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_95_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06846_ _01250_ _01288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_55_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09565_ net90 net8 _03729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06777_ _01218_ _01219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09638__A1 _03762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10248__A2 _04387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08516_ _02788_ _02789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_145_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09496_ _02809_ _00694_ _03663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_149_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_180_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08447_ as2650.stack\[15\]\[14\] _02706_ _02721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_24_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06872__A1 _01309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08378_ _02663_ _02667_ _02668_ _02671_ _00164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_139_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07329_ _01764_ _01765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08613__A2 _01195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09810__A1 _02094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06624__A1 _01063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10340_ _00737_ _02614_ _04343_ _04465_ _04456_ _04466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__10420__A2 _02570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10271_ _04409_ _03685_ _04307_ _04410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_84_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12010_ _00379_ clknet_leaf_117_wb_clk_i as2650.stack\[9\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_191_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10184__A1 _00801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_47_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10723__A3 _04831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09316__I _02626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_48_wb_clk_i clknet_4_13_0_wb_clk_i clknet_leaf_48_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_11725_ _00108_ clknet_leaf_86_wb_clk_i as2650.stack\[0\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08852__A2 _03067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06863__A1 _00709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11656_ _00039_ clknet_leaf_122_wb_clk_i as2650.stack\[11\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_70_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11721__CLK clknet_leaf_5_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout90 net55 net90 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_128_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10607_ _02619_ _04702_ _04717_ _04606_ _04718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_156_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09801__A1 _02859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11587_ _02101_ _05624_ _05631_ _05076_ _00413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__09801__B2 _03960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10538_ _04649_ _04650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_157_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_170_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11871__CLK clknet_leaf_38_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10469_ _04581_ _04582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_124_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08368__A1 _02527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07040__A1 _01478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06394__A3 _00667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08130__I _02466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09868__A1 _01609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06700_ _00930_ _00649_ _01143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_38_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09670__B _03832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10478__A2 _03866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07680_ as2650.stack\[13\]\[5\] _02025_ _02103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_65_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06631_ _01060_ _01074_ _01075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_1514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06585__I _05730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09350_ _02045_ _03548_ _02659_ _03549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__11427__A1 _03571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06562_ _01005_ _00634_ _00957_ _01006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08301_ net75 _02610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_21_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09281_ _03495_ _03496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_61_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06493_ _00936_ _00937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08232_ _02521_ _02541_ _02542_ _02543_ _00146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_60_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05901__I0 as2650.r123\[1\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08163_ _02492_ _02493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10835__I _02557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07114_ _01547_ _01551_ _01552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_140_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08305__I _02613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10402__A2 _02556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08094_ _02388_ _02437_ _02438_ _02439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_161_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06082__A2 as2650.cycle\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07045_ _01478_ _01481_ _01483_ _01484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_161_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08359__A1 as2650.stack\[3\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10166__A1 _03870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06909__A2 _01326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07031__A1 _01460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_5718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_173_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_130_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08996_ _03231_ _03222_ _03225_ _03232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_125_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07582__A2 _00929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07947_ _02213_ _02321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_131_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09859__A1 _04008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11115__B1 _05153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07878_ _02268_ _02269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_84_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08531__A1 _02793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07334__A2 _01769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09617_ _03654_ _03781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_56_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06829_ net10 _01271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_186_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11418__A1 _03561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09548_ _00703_ _01712_ _02580_ _03712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_77_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11744__CLK clknet_leaf_114_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_184_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_169_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09479_ _00541_ _03646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_93_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11433__A4 _01292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11510_ _01986_ _05165_ _05559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_169_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11441_ _05506_ _05507_ _00391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_138_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_109_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08598__A1 _02805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08215__I _02530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11372_ _02030_ _02137_ _02664_ _05455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_125_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10323_ _04452_ as2650.holding_reg\[7\] _04425_ _04453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_109_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10254_ _00978_ _04392_ _04398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_152_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09011__A2 _03233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10185_ _02893_ _04325_ _04335_ _00507_ _04336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_121_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08770__A1 _02388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10172__A4 _03695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05887__A2 _05740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11409__A1 as2650.stack\[9\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10880__A2 _04975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11244__C _05215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_15_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08825__A2 _00983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06836__A1 _01277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11708_ _00091_ clknet_leaf_127_wb_clk_i as2650.stack\[14\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_42_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10632__A2 _04703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09649__C _00552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11260__B _02814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11639_ _00022_ clknet_leaf_37_wb_clk_i as2650.r123\[0\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_128_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08589__A1 _02860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10396__A1 net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_32_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09250__A2 _02234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07261__A1 _05796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07964__I _02008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10148__A1 _02225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10604__B _04610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08850_ _01097_ _03096_ _03097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_48_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07801_ net66 _02211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08761__A1 _02412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08781_ _02368_ _03029_ _03034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_152_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05993_ _00451_ _00452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_113_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07732_ _02131_ _01729_ _02152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_66_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11767__CLK clknet_leaf_92_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08513__A1 as2650.stack\[5\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08513__B2 as2650.stack\[4\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07663_ _02036_ _02087_ _02063_ _02088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_81_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_187_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09402_ _02511_ _03589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06614_ _00652_ _01058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_25_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09069__A2 _03292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11154__C _05241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07594_ _05676_ _02018_ _02021_ _02022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_41_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09333_ _03040_ _03533_ _03534_ _03535_ _00255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_59_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06545_ _00988_ _00989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_107_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09264_ _03467_ _03469_ _03481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11281__C1 as2650.stack\[10\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06476_ net28 net15 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_139_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08292__A3 _02598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08215_ _02530_ _02531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_138_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09195_ _05759_ _03393_ _03415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08146_ _02323_ _02468_ _02474_ _02479_ _00124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__08035__I _02050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10387__A1 net47 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07252__A1 _01451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08077_ _02418_ _02427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_150_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07028_ _01466_ _00933_ _01467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_192_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11336__B1 _05154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07004__A1 _01316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07004__B2 _01318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_88_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_102_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06358__A3 _00646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08979_ _02648_ _02000_ _03218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_75_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11990_ _00359_ clknet_leaf_26_wb_clk_i as2650.r0\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_4869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_99_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10941_ _04916_ _05028_ _05042_ _03816_ _05043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_28_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10311__A1 _04327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10872_ _04199_ _04102_ _04676_ _04976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06818__A1 _00423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06953__I _05760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11272__C1 as2650.stack\[6\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09480__A2 _02759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07491__B2 as2650.stack\[13\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_8_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09768__B1 _03916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11424_ _03568_ _05487_ _05492_ _05493_ _00388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_184_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10378__A1 net45 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_177_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06046__A2 _00504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11355_ _05446_ _00366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_180_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10306_ _01905_ _04439_ _04440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_141_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11286_ _05189_ _05363_ _05379_ _05380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_10237_ _02845_ _04157_ _04385_ _04386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_140_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10168_ _00556_ _00715_ _03650_ _04319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_94_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10550__A1 _00780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10099_ _04249_ _04251_ _04252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__09299__A2 _03502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_63_wb_clk_i clknet_4_15_0_wb_clk_i clknet_leaf_63_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_130_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07959__I _02236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06330_ _00779_ _00780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_188_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06261_ _00712_ _00625_ _00715_ _00716_ _00001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_31_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08000_ _02364_ _02365_ _02366_ _02367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_102_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06192_ _05728_ _00651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09223__A2 _01518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07694__I _02115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08982__A1 as2650.stack\[7\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09951_ _02126_ _04101_ _04107_ _04108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_143_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11318__B1 _05401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08902_ _03110_ _03145_ _03146_ _00213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09882_ _04024_ _04032_ _04033_ _04039_ _04040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_135_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08734__A1 _02003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08833_ _03079_ _03080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_22_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08739__B _02701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10988__C _04904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_170_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08764_ _02415_ _03011_ _03018_ _03019_ _00202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05976_ _05791_ _00434_ _00431_ _00435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_57_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07715_ _02134_ _02135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11097__A2 _05194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08695_ _02925_ _02966_ _02967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_38_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_148_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07646_ _01263_ _02042_ _02072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__10844__A2 net88 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07577_ _00554_ _00904_ _02005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_126_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09316_ _02626_ _03523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_90_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_139_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06528_ _00694_ _00971_ _00972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_40_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_194_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09462__A2 _03627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07473__A1 _01905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09247_ _03393_ _03465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06459_ _00645_ _00904_ _00905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08670__B1 _01435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_194_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_177_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_166_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09178_ _03397_ _03398_ _03399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_147_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11557__B1 _05601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08129_ _02465_ _02249_ _02466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07076__I1 as2650.r123_2\[0\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11021__A2 _04309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08973__A1 _01693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput23 net23 io_out[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_190_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11140_ _04275_ _01261_ _05237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_122_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput34 net34 io_out[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_150_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11932__CLK clknet_leaf_61_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xoutput45 net45 io_out[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__10780__A1 _03921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11309__B1 _05172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput56 net56 la_data_out[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_122_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput67 net67 la_data_out[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_89_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput78 net78 la_data_out[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_11071_ _05151_ _05170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_5301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output65_I net87 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08725__A1 _02409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_172_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10022_ _04175_ _04176_ _04177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__08725__B2 _02990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_193_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_102_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06200__A2 _00505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11973_ _00342_ clknet_leaf_50_wb_clk_i net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_4688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10924_ _05025_ _05026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_44_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10855_ _04952_ _04954_ _04959_ _04960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_44_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__10599__A1 _03921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10786_ _04883_ _04885_ _04887_ _04892_ _04893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_12_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09453__A2 _03615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_140_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07464__B2 as2650.stack\[8\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06019__A2 _00477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11407_ _02364_ _05480_ _05481_ _05482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__11012__A2 _00973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08964__A1 as2650.r123_2\[1\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10220__B1 _04360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08403__I _02689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11338_ _05428_ _05429_ _05430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11563__A3 _02734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_4_9_0_wb_clk_i clknet_3_4_0_wb_clk_i clknet_4_9_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_67_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_154_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09943__B _03728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11269_ _05351_ _05362_ _02805_ _05363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_171_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_84_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07019__I _01457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07519__A2 _01832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08716__A1 _02452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10523__A1 _01765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05830_ _05683_ _05684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_23_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07463__B _01846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05950__A1 _05802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07500_ as2650.r123\[0\]\[5\] _01931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_149_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10826__A2 _04931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08480_ _00831_ _00768_ _02753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09692__A2 _03852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07431_ _01824_ _01865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_126_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11805__CLK clknet_leaf_3_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07362_ _01783_ _01785_ _01797_ _01798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_189_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09444__A2 _03613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08247__A3 _00658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09101_ _05764_ _01515_ _03324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_148_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06313_ _00656_ _00764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_149_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06258__A2 _00713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08652__B1 _02923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07293_ net48 _01729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11251__A2 _05345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_191_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_176_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09032_ _03249_ _03262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06244_ _00492_ _00457_ _00701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_190_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11955__CLK clknet_leaf_20_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07207__A1 as2650.r0\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10843__I _03665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06175_ as2650.cycle\[9\] _00632_ _00634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10762__B2 _04534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09934_ _00719_ _04086_ _04090_ _03777_ _04091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA_clkbuf_leaf_59_wb_clk_i_I clknet_4_15_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08707__A1 _02976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09865_ _02115_ _04023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10514__A1 as2650.stack\[1\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10514__B2 as2650.stack\[0\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09380__A1 as2650.stack\[3\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08816_ _03062_ _03063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09796_ _00717_ _03936_ _03955_ _02890_ _03956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__06194__A1 as2650.ins_reg\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06733__A3 _01173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08747_ _02449_ _03001_ _03005_ _03008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05959_ _05807_ _05812_ _05813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_45_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08678_ _02926_ _02936_ _02937_ _02949_ _02950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__10817__A2 _04922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09683__A2 _03844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07629_ _02055_ _02056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07599__I _01771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10640_ _02093_ _04704_ _04750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_167_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06249__A2 _00705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08643__B1 _02914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10571_ as2650.stack\[5\]\[2\] _02913_ _02914_ as2650.stack\[4\]\[2\] _04683_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__11242__A2 _05336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08643__C2 _02799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_154_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06008__I net72 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11996__D _00365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09199__A1 _05731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_98_wb_clk_i_I clknet_4_9_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10753__A1 _00780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_194_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11123_ _00823_ _05221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_174_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06421__A2 _00763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11054_ _01855_ _05153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_5131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06709__B1 _01149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10505__A1 _04609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10005_ _03661_ _04161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_188_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06678__I _01009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06185__A1 _00625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11828__CLK clknet_leaf_34_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09989__I _02889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08893__I _01034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11956_ _00325_ clknet_leaf_17_wb_clk_i as2650.holding_reg\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_33_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08477__A3 _00616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10907_ _04596_ _05009_ _05010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07685__A1 _01954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11533__B _05192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11887_ _00256_ clknet_leaf_103_wb_clk_i as2650.stack\[4\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_177_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11252__C _05278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10838_ _03972_ _04943_ _04944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_13_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11233__A2 _02867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09938__B _02890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10769_ _02115_ _04007_ _04791_ _04876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_125_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10992__A1 _04439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08937__A1 _02836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06948__B1 _01387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10744__A1 _00894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08401__A3 _02664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07980_ _02348_ _02349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07972__I _00476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06931_ _00999_ _01351_ _01371_ _00017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_110_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08165__A2 _02489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09650_ _02889_ _03813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06862_ _01302_ _01303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_67_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06176__A1 _00511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08601_ _01660_ _01661_ _02874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_67_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07912__A2 _02297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09581_ _01130_ _03745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_83_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06793_ as2650.holding_reg\[2\] _00655_ _01232_ _01235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
Xwrapped_as2650_108 io_oeb[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_110_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08532_ _02777_ _02805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xwrapped_as2650_119 io_out[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_24_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09665__A2 _03752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07676__A1 _02091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08463_ _02731_ _02734_ _02735_ _02736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__11472__A2 _05531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_184_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07414_ _01801_ _01849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_51_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08394_ _02680_ _02681_ _02682_ _02683_ _00168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_52_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_132_wb_clk_i_I clknet_4_0_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09417__A2 _03599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07212__I _01648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07345_ _01780_ _01781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_91_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11224__A2 _01429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10432__B1 _02794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07276_ _00605_ _01711_ _01712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_191_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_163_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10983__A1 _00622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09015_ _00848_ _03101_ _03246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_152_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06227_ _00448_ _05680_ _00685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_164_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08928__A1 _01445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06158_ _00613_ _00616_ _00508_ _00617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_144_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10735__A1 _04007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06089_ _00536_ _00548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09917_ _04071_ _04072_ _04073_ _04074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_132_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09353__A1 _02284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11337__C _05364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09848_ net61 _04007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_115_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07364__B1 _01798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_160_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09779_ _03937_ _03938_ _03939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_27_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09105__A1 _05731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11810_ _00193_ clknet_leaf_5_wb_clk_i as2650.stack\[15\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09602__I _00991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output28_I net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11741_ _00124_ clknet_leaf_116_wb_clk_i as2650.stack\[8\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11463__A2 _05672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_187_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_148_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11672_ _00055_ clknet_leaf_131_wb_clk_i as2650.stack\[13\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_42_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08218__I _02533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09408__A2 _03589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10623_ _04732_ _04733_ _01776_ _04734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_139_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11215__A2 _05226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10423__B1 _01744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10554_ _04432_ _04661_ _04374_ _04666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_167_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10974__A1 _04532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10483__I _04595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10974__B2 _03757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07278__B _01052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10485_ _02057_ _02039_ _00804_ _04598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_5_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_170_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10726__A1 _02906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09592__A1 _03728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08888__I _03077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11106_ _05200_ _01195_ _05201_ _05203_ _05204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_61_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11650__CLK clknet_leaf_134_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11037_ _05135_ _04553_ _05136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06158__A1 _00613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_168_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08837__B _03079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__12006__CLK clknet_leaf_117_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_181_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11939_ _00308_ clknet_leaf_66_wb_clk_i net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_146_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07130_ as2650.holding_reg\[6\] _01568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_146_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_173_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10965__A1 _02229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07061_ _01059_ _01496_ _01499_ _01500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__06633__A2 _00515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07830__A1 _02234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07830__B2 _02235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06012_ _00466_ _00470_ _00471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_161_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10717__A1 as2650.stack\[3\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10717__B2 as2650.stack\[0\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08386__A2 _02667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09583__A1 _03732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08798__I _02112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07963_ _02331_ _02332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_141_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08138__A2 _02468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09335__A1 _02989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_190_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06914_ _01328_ _05752_ _01110_ _01212_ _01355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_09702_ _03729_ _03862_ _03863_ _03864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_116_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07894_ _02059_ _02284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__11142__A1 _05238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09886__A2 _04043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09633_ _03795_ _03796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_06845_ _01133_ _01286_ _01287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07897__A1 _02284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10996__C _04744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09564_ _03727_ _03728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06776_ _01217_ _01218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_55_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08515_ _02134_ _01736_ _02788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_164_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11445__A2 _03431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09495_ _03661_ _03662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_164_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08446_ _02684_ _02717_ _02718_ _02720_ _00183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_51_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08038__I _02256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08377_ _02670_ _02671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07328_ _01732_ _01764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_164_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_164_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08613__A3 _01249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09810__A2 _03725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07259_ _01695_ _01696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07821__A1 _02222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10270_ _03991_ _04409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_151_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10708__A1 _00522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09574__A1 _03723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11673__CLK clknet_leaf_131_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10184__A2 _04329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08129__A2 _02249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09326__A1 _03033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11067__C _05165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11133__A1 _05177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12029__CLK clknet_4_4_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09877__A2 _01473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10892__B1 _04979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_185_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06560__A1 _00540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05860__I _05713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11724_ _00107_ clknet_leaf_113_wb_clk_i as2650.stack\[0\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_175_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11655_ _00038_ clknet_leaf_126_wb_clk_i as2650.stack\[11\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06863__A2 _00585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout80 net82 net80 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_128_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout91 net27 net91 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06691__I _05781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10606_ _05673_ _04711_ _04717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_88_wb_clk_i clknet_4_8_0_wb_clk_i clknet_leaf_88_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__08065__A1 _02415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11586_ _05413_ _04837_ _05624_ _05630_ _05631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_10_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09801__A2 _03872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06624__C _01067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_17_wb_clk_i clknet_4_5_0_wb_clk_i clknet_leaf_17_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_10537_ _04648_ _04649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10411__A3 _04341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11102__I _00774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10468_ _02056_ _03722_ _04581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_174_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_170_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09565__A1 net90 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10399_ _02347_ _04483_ _04513_ _04514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_97_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11372__A1 _02030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07040__A2 _00830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09317__A1 _03000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09868__A2 _01618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07027__I _01465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06630_ _01069_ _01073_ _01074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06866__I _01027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06561_ _00722_ _01004_ _01005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10388__I _04404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11427__A2 _05487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08300_ _01459_ _02608_ _02609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_61_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09280_ _02272_ _02437_ _03024_ _03495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_06492_ _00746_ _00469_ _00936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_94_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08231_ as2650.stack\[5\]\[12\] _02538_ _02543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__06854__A2 _01295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05901__I1 as2650.r123\[0\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07697__I _02118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08162_ _02133_ _02491_ _02471_ _02492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__08056__A1 _02177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10938__A1 _02216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07113_ _01548_ _01549_ _01550_ _01551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_88_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08093_ _02022_ _02438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07803__A1 _01219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07803__B2 _02212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10402__A3 _03702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07044_ _05740_ _00991_ _01482_ _00656_ _01483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__08359__A2 _02655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10166__A2 _00812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_173_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08995_ _02086_ _03231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_29_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09308__A1 _02184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07946_ _02318_ _02315_ _02320_ _02317_ _00083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_5_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06790__A1 _00421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11115__A1 as2650.stack\[6\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11115__B2 as2650.stack\[5\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07877_ _02198_ _02136_ _02254_ _02268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__06917__I0 as2650.r123\[0\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08531__A2 _02803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09616_ _03779_ _03780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06828_ _00426_ _01045_ _01270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_28_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11615__C _00712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06709__C _00943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06759_ _01135_ _01021_ _01111_ _01201_ _01202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__11418__A2 _05487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09547_ _03710_ _03711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_43_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10626__B1 _01780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08991__I _03219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_180_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09478_ _00564_ _03644_ _03645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_54_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06845__A2 _01286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08429_ _02133_ _02491_ _01995_ _02709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
Xclkbuf_4_11_0_wb_clk_i clknet_3_5_0_wb_clk_i clknet_4_11_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_106_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11440_ _01808_ _05499_ _05504_ as2650.r123\[2\]\[1\] _05507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08047__A1 _02170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07400__I _01809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09795__A1 _03759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11371_ _05454_ _00374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09795__B2 _03772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10322_ _02903_ _00795_ _02353_ _04452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_180_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07270__A2 _01686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10253_ _02933_ _04397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_140_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_191_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11354__A1 _02625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05855__I net51 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07022__A2 _05748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10184_ _00801_ _04329_ _04330_ _04334_ _04335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_61_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08770__A2 _02146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_135_wb_clk_i clknet_4_1_0_wb_clk_i clknet_leaf_135_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_19_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11409__A2 _05478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_182_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10001__I _04156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08286__A1 _00597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08825__A3 _03054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_148_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10093__A1 _04209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11707_ _00090_ clknet_leaf_127_wb_clk_i as2650.stack\[14\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11638_ _00021_ clknet_leaf_35_wb_clk_i as2650.r123\[1\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_129_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11260__C _00842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07310__I _01745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09786__A1 _03165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08589__A2 _02613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11569_ _01675_ _05614_ _05615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_6_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09538__A1 _00467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11345__A1 _05364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09553__A4 _03716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07800_ _02189_ _02207_ _02209_ _02210_ _00047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__08761__A2 _03011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08780_ _02066_ _03033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_85_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_111_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05992_ _00450_ _00451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_111_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07980__I _02348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07731_ _02044_ _02151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_78_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08513__A2 _02785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07662_ _02086_ _02087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_113_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06524__A1 _00955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06613_ _01007_ _01012_ _01056_ _01057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09401_ _03558_ _03575_ _03587_ _03588_ _00270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_65_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07593_ _02019_ _02020_ _02021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_74_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06544_ as2650.idx_ctrl\[1\] as2650.idx_ctrl\[0\] _00988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_09332_ _02456_ _03523_ _03527_ _03535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_181_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10084__A1 _02212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09263_ _02345_ _03465_ _03440_ _03480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__10084__B2 _04237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11281__B1 _01914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06475_ _00452_ _00821_ _00890_ _05674_ _00920_ _00000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_37_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11281__C2 _01912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08214_ _02529_ _02530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_53_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09194_ _03412_ _03413_ _03414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_166_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09777__A1 _02853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08145_ as2650.stack\[8\]\[11\] _02477_ _02479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_135_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11584__A1 _01462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08076_ _02318_ _02420_ _02424_ _02426_ _00107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_161_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09529__A1 _02599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07027_ _01465_ _01466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_118_1511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11336__A1 as2650.stack\[5\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11336__B2 as2650.stack\[7\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_161_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07004__A2 _01424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08201__A1 _02519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_142_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09544__A4 _03672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_5538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06763__A1 _01202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08978_ _03216_ _03217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_76_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_102_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07890__I _02280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_102_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11626__B _02340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07929_ _02304_ _02214_ _02309_ _02306_ _00077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_4859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10940_ _04806_ _05041_ _05042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06515__A1 _00772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10311__A2 _04394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08000__B _02366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10871_ _04223_ _04974_ _04975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_45_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08268__A1 _02012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09610__I _00551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__11272__B1 _05303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__11272__C2 _05296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_185_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07491__A2 _01874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07130__I as2650.holding_reg\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09768__A1 _03914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11423_ _02119_ _05462_ _05472_ _05493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_172_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11575__A1 _04161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11354_ _02625_ _05444_ _05445_ _05446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__07243__A2 _01583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08440__A1 _02678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10705__B _04105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10305_ _04428_ _04439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_119_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10491__I _02824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11285_ _05152_ _05370_ _05378_ _05185_ _05379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_153_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11327__A1 _02951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10236_ _04384_ _04385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_3_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_171_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10167_ _00891_ _04317_ _03598_ _04318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_67_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10550__A2 _04648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10098_ _04250_ _04218_ _04251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_3_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10302__A2 _04435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_130_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07305__I net86 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_169_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10066__A1 _00633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11271__B _05364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_32_wb_clk_i clknet_4_7_0_wb_clk_i clknet_leaf_32_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_124_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06260_ _00530_ _00692_ _00716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06191_ _00649_ _00612_ _00650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_11_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09950_ _04102_ _04089_ _04106_ _04107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_104_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11318__A1 _00824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08901_ _01222_ _03108_ _03130_ as2650.r123_2\[1\]\[2\] _03146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_clkbuf_leaf_49_wb_clk_i_I clknet_4_13_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09881_ _03894_ _04038_ _03794_ _04039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09931__A1 net36 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08832_ _01143_ _03076_ _03079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10541__A2 _04597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05975_ _05809_ _00434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08763_ _02302_ _02695_ _02995_ _03019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_73_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10350__B _00467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07714_ net70 _02134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_66_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08498__A1 _02747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08694_ _02843_ _02963_ _02965_ _02966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_26_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07645_ _02070_ _02071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_26_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07576_ _00925_ _02004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_40_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10057__A1 _04209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06527_ _00561_ _00971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__09998__A1 _04131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09315_ as2650.stack\[4\]\[0\] _03521_ _03522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_139_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09246_ _03461_ _03463_ _03464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_139_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06458_ as2650.cycle\[4\] _00561_ _00904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__08670__A1 _02065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08670__B2 _02089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09177_ _05732_ _01517_ _03398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_88_wb_clk_i_I clknet_4_8_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06389_ _00834_ _00835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11557__A1 _00754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07885__I _02044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08128_ _01933_ _02145_ _02465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11557__B2 _02740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08422__A1 _02684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput13 net13 io_oeb[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_08059_ as2650.stack\[12\]\[6\] _02396_ _02413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xoutput24 net24 io_out[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_85_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput35 net35 io_out[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_159_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11200__I _01862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11309__A1 as2650.stack\[9\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput46 net46 io_out[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__06984__A1 _01390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11309__B2 as2650.stack\[11\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10780__A2 _00895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput57 net89 la_data_out[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11070_ _05155_ _05161_ _05168_ _05169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xoutput68 net68 la_data_out[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_163_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput79 net79 la_data_out[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_5302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_5313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10021_ _04156_ _04124_ _04126_ _04176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_103_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09922__A1 _04078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08725__A2 _02985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output58_I net58 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06200__A3 _00614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08489__A1 _00754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11972_ _00341_ clknet_leaf_39_wb_clk_i net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_4689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11088__A3 _05186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_99_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10923_ _02224_ _05025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_3988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10854_ _04590_ _04956_ _04958_ _04891_ _04959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_16_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_144_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_164_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10785_ _04808_ _04889_ _04890_ _04891_ _04892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_38_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10599__A2 _03920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_73_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_157_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_157_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07464__A2 _01869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11548__A1 _05589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11548__B2 _04298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11757__CLK clknet_leaf_80_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11406_ _05460_ _05481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07216__A2 _01652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08413__A1 as2650.stack\[1\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11012__A3 _00986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10220__A1 _00707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11337_ as2650.stack\[6\]\[7\] _05212_ _05157_ as2650.stack\[4\]\[7\] _05364_ _05429_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__11563__A4 _05608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06975__A1 _01086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_193_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06975__B2 _01088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06204__I _00589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11268_ _01463_ _00789_ _05205_ _02835_ _05361_ _05362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_49_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09913__A1 _01610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08716__A2 _02974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10219_ _04366_ _04368_ _04349_ _04369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_11199_ as2650.stack\[5\]\[3\] _05162_ _05163_ as2650.stack\[7\]\[3\] _05295_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_132_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11266__B _05359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07035__I _01473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07152__A1 _05802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07430_ as2650.stack\[3\]\[10\] _01862_ _01863_ as2650.stack\[0\]\[10\] _01753_ as2650.stack\[1\]\[10\]
+ _01864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_23_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_22_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10039__A1 _04109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_122_wb_clk_i_I clknet_4_0_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07361_ _01788_ _01792_ _01796_ _01797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_17_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11236__B1 _05163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09100_ as2650.r0\[2\] _01542_ _03323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06312_ _00479_ _00763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08247__A4 _02555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07292_ _01727_ _01728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_148_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08652__A1 _02912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_148_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08652__B2 _01845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09031_ _01203_ _03261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06243_ _00520_ _00699_ _00700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07919__B _02269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_1811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_1822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_1833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07207__A2 _01358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06174_ _00632_ _00633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__11003__A3 _03686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_5_wb_clk_i_I clknet_4_1_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10211__A1 _04331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_1888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10762__A2 _02804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09933_ _03772_ _04089_ _04090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_131_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08707__A2 _02717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09864_ _03974_ _04022_ _00299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_112_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_154_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10514__A2 _01829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08815_ _01129_ _01131_ _03061_ _03062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XTAP_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09795_ _03759_ _03950_ _03954_ _03772_ _03789_ _03955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XTAP_3207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_96_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08746_ as2650.stack\[1\]\[2\] _02998_ _03007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05958_ _05808_ _05770_ _05785_ _05810_ _05811_ _05812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_113_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05941__A2 _05749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10278__A1 _02865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05889_ _05742_ _05743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07143__A1 _01480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08677_ _02938_ _02943_ _02926_ _02948_ _02949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06784__I _00968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07628_ _02054_ _02055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_26_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08891__A1 _02849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07559_ _00605_ _00974_ _01986_ _01987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_195_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_167_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10570_ as2650.stack\[7\]\[2\] _02799_ _04681_ as2650.stack\[6\]\[2\] _04682_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_107_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07446__A2 _01816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08643__A1 as2650.stack\[1\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08643__B2 as2650.stack\[0\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_155_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09229_ _03424_ _03448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_194_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_166_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_155_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09199__A2 _02233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08504__I _00865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_182_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10202__A1 _03710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06957__A1 _01392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10753__A2 _04859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11122_ _05214_ _05219_ _05152_ _05220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_122_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06421__A3 _00849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11053_ _05151_ _05152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_77_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06709__A1 _01139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10505__A2 _04582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10004_ _02195_ _03959_ _04159_ _03968_ _04160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_5154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_123_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09123__A2 _03333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10269__A1 _03712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11955_ _00324_ clknet_leaf_20_wb_clk_i as2650.holding_reg\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08477__A4 _01130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06694__I _00943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10906_ _04999_ _05008_ _05009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_32_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08882__A1 _01195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06488__A3 _00927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11533__C _02350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11886_ _00255_ clknet_leaf_98_wb_clk_i as2650.stack\[4\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_33_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10837_ _04937_ _04940_ _04942_ _04943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_60_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_157_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07437__A2 _01869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10768_ net63 _04875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__10441__A1 _03722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07739__B _02158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10699_ _00779_ _04808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_195_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06948__B2 _01223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09673__C _03786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_190_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06930_ as2650.r123\[1\]\[3\] _01197_ _01370_ _01207_ _01371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_141_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06869__I net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input1_I io_in[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06861_ _01297_ _01010_ _01298_ _01299_ _01300_ _01301_ _01302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_67_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06176__A2 _00630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08600_ _01572_ _01678_ _02873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_27_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06792_ _01227_ _01234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09580_ _03743_ _03744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_95_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_110_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xwrapped_as2650_109 io_oeb[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_188_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08531_ _02793_ _02803_ _02804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_149_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08462_ _00773_ _00964_ _00982_ _02735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_23_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07676__A2 _02092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11922__CLK clknet_leaf_49_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07413_ _01203_ _01803_ _01848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_50_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08393_ as2650.stack\[2\]\[12\] _02676_ _02683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_50_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07344_ _01779_ _01780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06109__I net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10432__A1 as2650.stack\[9\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07275_ _05681_ _05670_ _01711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10432__B2 as2650.stack\[8\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07649__B _02063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09014_ _03244_ _03245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06226_ _00678_ _00680_ _00683_ _00684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__10983__A2 _00699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08324__I _02631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06157_ _00615_ _00616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_195_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_191_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06088_ _00541_ _00546_ _00547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_78_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09916_ _04071_ _04072_ _03887_ _04073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_115_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11618__C _05658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09847_ _03977_ _02890_ _04005_ _04006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XTAP_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09778_ _02852_ _01302_ _03842_ _03843_ _03889_ _03938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XTAP_3026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09105__A2 _01358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08729_ _02381_ _02974_ _02993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07116__B2 _01357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11740_ _00123_ clknet_leaf_116_wb_clk_i as2650.stack\[8\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10671__A1 as2650.stack\[11\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11671_ _00054_ clknet_leaf_130_wb_clk_i as2650.stack\[13\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_14_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10622_ as2650.stack\[3\]\[3\] _01839_ _02907_ _04733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_128_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_155_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10423__A1 as2650.stack\[7\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10423__B2 as2650.stack\[6\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10553_ _04652_ _04657_ _04664_ _04665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_10_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10484_ net90 as2650.ins_reg\[2\] net56 _04597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_183_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09041__A1 _03145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_139_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09493__C _03659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11105_ _03948_ _01161_ _05202_ _05203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_1_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11036_ _00847_ _05135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06158__A2 _00616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11945__CLK clknet_leaf_54_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07107__A1 _05781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_146_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11938_ _00307_ clknet_leaf_38_wb_clk_i net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08855__A1 _00835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08409__I _02688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10662__A1 _04609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11869_ _00238_ clknet_leaf_34_wb_clk_i as2650.r123_2\[2\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_18_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_158_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09280__A1 _02272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10965__A2 _05064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07060_ _01341_ _01497_ _01489_ _01498_ _01166_ _01499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__10607__C _04606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_103_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06011_ _00469_ _00470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_173_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05841__A1 _05691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_160_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09684__B _01002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07983__I _02351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10717__A2 _04822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10623__B _01776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07594__A1 _05676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06599__I _01042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07962_ _05671_ _02331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09701_ _02054_ _03790_ _03863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06913_ _01328_ _01110_ _01212_ _05814_ _01354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_9_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09335__A2 _02634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07893_ as2650.stack\[10\]\[1\] _02274_ _02283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11142__A2 _01286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09632_ net9 _03795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_95_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06844_ _01281_ _01283_ _01285_ _01286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_83_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_83_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09563_ _00804_ _02865_ _00816_ _03727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_110_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06775_ _01216_ _01217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_110_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08514_ _01733_ _02783_ _02786_ _02787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_70_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11173__C _05215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08319__I _02626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07649__A2 _02074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09494_ _02807_ _03661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_145_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10653__A1 _02852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08445_ as2650.stack\[15\]\[13\] _02714_ _02720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_145_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08376_ _02669_ _02670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10405__A1 _04351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07327_ as2650.stack\[3\]\[8\] _01740_ _01761_ as2650.stack\[0\]\[8\] _01762_ as2650.stack\[1\]\[8\]
+ _01763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XANTENNA__09271__A1 _02346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08613__A4 _01350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08054__I _02101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07258_ _01601_ _01017_ _01688_ _01319_ _01694_ _01695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_10_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07821__A2 _02227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05832__A1 _05682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06209_ _00651_ _00667_ _00668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11818__CLK clknet_4_3_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07189_ _01533_ _01624_ _01625_ _01626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09023__A1 _01101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09594__B _03756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07034__B1 _01456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09574__A2 _05672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07826__C _02201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07585__A1 _00948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06730__C _01067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11381__A2 _05462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07337__A1 _01771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_output40_I net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09613__I _03776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10892__A1 _01884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10892__B2 _03667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06560__A2 _00720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08837__A1 _00428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08229__I _02530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10644__A1 _03921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11723_ _00106_ clknet_leaf_83_wb_clk_i as2650.stack\[0\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09769__B _03883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06972__I _01396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11654_ _00037_ clknet_leaf_3_wb_clk_i as2650.stack\[13\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06863__A3 _00642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout81 net82 net81 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_174_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout92 net42 net92 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_10605_ _04584_ _04707_ _04713_ _04715_ _04716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_155_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08065__A2 _02406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11585_ _05553_ _05625_ _05629_ _00756_ _05630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_7_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10536_ _04646_ _04647_ _04648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_176_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07812__A2 _02208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_155_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10467_ _03726_ _04531_ _04580_ _04506_ _00344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_124_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09565__A2 net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11539__B _04501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_57_wb_clk_i clknet_4_15_0_wb_clk_i clknet_leaf_57_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_151_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10398_ _02834_ _04484_ _04513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_124_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10580__B1 _02914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09317__A2 _03523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11019_ _05117_ _05118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_113_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06551__A2 _00975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06560_ _00540_ _00720_ _01004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08139__I _02466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10635__A1 _02082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06491_ _00479_ _00872_ _00935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_61_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07978__I _02346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08230_ _02534_ _02542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_166_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05901__I2 as2650.r123_2\[1\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10650__A4 _04759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08161_ _01988_ _02491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_147_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08056__A2 _02258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07112_ _05765_ _01359_ _01550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08092_ _01769_ _02437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_147_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_146_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07043_ _05733_ _00962_ _01482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09005__A1 as2650.stack\[7\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10166__A3 _03651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_134_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08994_ as2650.stack\[7\]\[3\] _03220_ _03230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10571__B1 _02914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09308__A2 _03502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07945_ as2650.stack\[10\]\[9\] _02319_ _02320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_130_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11115__A2 _05212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07876_ _02237_ _02263_ _02264_ _02267_ _00066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_44_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09615_ _00730_ _03779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06827_ _01268_ _01269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_112_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10874__A1 _04223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06542__A2 _00631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08049__I _02090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09546_ _03707_ _03709_ _03710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06758_ _01200_ _01201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08819__A1 _00987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10626__A1 as2650.stack\[15\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10626__B2 as2650.stack\[14\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09477_ _00928_ _00772_ _03644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09589__B _03723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08295__A2 _02590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06689_ _00942_ _01129_ _01131_ _01132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__09492__A1 _02568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07888__I _02278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06792__I _01227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08428_ as2650.stack\[15\]\[8\] _02706_ _02708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_157_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10528__B _04639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11640__CLK clknet_leaf_36_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08359_ as2650.stack\[3\]\[11\] _02655_ _02657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08047__A2 _02392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10929__A2 _02216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06058__A1 _00449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07255__B1 _01688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11051__A1 _01992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11370_ as2650.r123_2\[3\]\[7\] _05454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09795__A2 _03950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10321_ _04451_ _00327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_193_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06741__B _01031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_49_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10252_ _04394_ _04387_ _04396_ _00313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08512__I _02784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10183_ net28 _04333_ _03968_ _04334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_152_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06032__I _05691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11106__A2 _01195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09343__I _01030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10865__A1 _04948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07730__A1 as2650.stack\[11\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_104_wb_clk_i clknet_4_3_0_wb_clk_i clknet_leaf_104_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_131_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08286__A2 _00603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11290__A1 _03761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11706_ _00089_ clknet_4_4_0_wb_clk_i net77 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07494__B1 _01925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_188_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_175_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11637_ _00020_ clknet_leaf_36_wb_clk_i as2650.r123\[1\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_180_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06049__A1 _00506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11042__A1 _02819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09786__A2 _01445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08589__A3 _02861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11568_ _01674_ _01672_ _05614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_7_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_171_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_155_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10519_ as2650.stack\[11\]\[1\] _01835_ _01823_ as2650.stack\[10\]\[1\] _04632_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_143_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11499_ _05551_ _00405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_100_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__11269__B _02805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_39_wb_clk_i_I clknet_4_6_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05991_ _00449_ _00450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_38_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07730_ as2650.stack\[11\]\[0\] _02149_ _02150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_133_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10856__A1 _04116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07661_ _02082_ _02083_ _02085_ _02086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_26_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06524__A2 _00957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09400_ _02087_ _02514_ _03582_ _03588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_65_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06612_ _01014_ _01019_ _01054_ _01055_ _01056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_25_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07592_ _00861_ _01104_ _02020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10608__A1 net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09331_ as2650.stack\[4\]\[4\] _03521_ _03534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06543_ _00985_ _00554_ _00986_ _00987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_94_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08277__A2 _02584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06288__A1 _00581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09262_ _03463_ _03478_ _03479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10084__A2 _04008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07485__B1 _01863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11281__A1 as2650.stack\[9\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06474_ _00556_ _00892_ _00918_ _00919_ _00920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_33_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11281__B2 as2650.stack\[8\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_194_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07501__I _01502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08213_ _02030_ _02485_ _02486_ _02529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_124_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09193_ _03392_ _03400_ _03413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09226__A1 _01663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08029__A2 _02001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_140_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11033__A1 net78 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09777__A2 _01302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08144_ _02321_ _02468_ _02474_ _02478_ _00123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_88_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11584__A2 _02833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08075_ as2650.stack\[0\]\[9\] _02425_ _02426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07252__A3 _01461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07026_ _01464_ _01465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09529__A2 _03691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11336__A2 _05153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09872__B _03766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05892__S _05713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06212__A1 _00662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08977_ _02492_ _03216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_4805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_2_wb_clk_i clknet_4_1_0_wb_clk_i clknet_leaf_2_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_4838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07928_ as2650.stack\[11\]\[10\] _02307_ _02309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_29_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09701__A2 _03790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07859_ _02256_ _02257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_57_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06515__A2 _00958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10870_ net65 net64 _04914_ _04974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_72_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_164_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09529_ _02599_ _03691_ _02549_ _03692_ _03693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_25_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08268__A2 _00841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09465__A1 _03568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06279__A1 _00707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11272__A1 as2650.stack\[5\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_101_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11272__B2 as2650.stack\[7\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07411__I _01845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_184_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09217__A1 _05733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_8_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11422_ as2650.stack\[9\]\[6\] _05476_ _05492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11024__A1 _02734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09768__A2 _03725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11575__A2 _05616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10772__I _00782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11353_ _02347_ _05148_ _05445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__08440__A2 _02707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_180_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06451__A1 _00686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10304_ _02332_ _04437_ _04438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_141_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11284_ _05170_ _05377_ _05378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11327__A2 _00874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09782__B _00534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10235_ _04372_ _04373_ _04383_ _04384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_106_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10166_ _03870_ _00812_ _03651_ _04311_ _04317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_94_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07951__A1 as2650.stack\[10\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05962__B1 _05755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10097_ _02211_ _04229_ _04250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_23_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09153__B1 _03374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10838__A1 _03972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11686__CLK clknet_leaf_124_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10012__I net87 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_112_wb_clk_i_I clknet_4_3_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10999_ _02841_ _02772_ _05097_ _00951_ _05098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_147_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__11263__A1 _05249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08417__I _02689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_187_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_176_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10605__A4 _04715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07321__I _01756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11015__A1 _00864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06190_ _00588_ _00593_ _00649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_72_wb_clk_i clknet_4_11_0_wb_clk_i clknet_leaf_72_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_102_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11566__A2 _01583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10615__C _04725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06442__A1 _00882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11318__A2 _05394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08900_ _03069_ _03143_ _03144_ _03145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_131_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09880_ _04034_ _04037_ _04038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_139_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_8_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08831_ _03077_ _03078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_97_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09931__A2 net35 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08734__A3 _02147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07924__C _02306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07942__A1 _02314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08762_ as2650.stack\[1\]\[7\] _03004_ _03018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05974_ _05791_ _00431_ _00432_ _00433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_39_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10829__A1 _05673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07713_ _02132_ _02133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_38_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09695__A1 _03836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08693_ _02964_ _02965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08498__A2 _02337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_26_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07644_ _02069_ _02070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_53_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07575_ _02002_ _02003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_53_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09314_ _03520_ _03521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06526_ _00946_ _00970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07458__B1 _01859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09998__A2 _03867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08327__I _02626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_178_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09245_ _03444_ _03462_ _03463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_178_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06457_ _00468_ _00550_ _00713_ _00530_ _00903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_107_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08670__A2 _02848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11006__A1 _00766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_193_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06681__A1 _01120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_182_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09176_ _03394_ _03396_ _03397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_06388_ _00658_ _00834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_120_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11557__A2 _04621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08127_ _02415_ _02454_ _02463_ _02464_ _00120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_179_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08422__A2 _02700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08062__I _02121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput14 net14 io_oeb[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_11_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08058_ _02112_ _02412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput25 net25 io_out[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_135_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput36 net36 io_out[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_134_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11309__A2 _05171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput47 net47 io_out[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_172_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07009_ _01226_ _01422_ _01448_ _01449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_116_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput58 net58 la_data_out[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_81_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput69 net69 la_data_out[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_131_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08186__A1 as2650.stack\[6\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10020_ _04174_ _04175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_5314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06736__A2 _01173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07933__A1 _02161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_5369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06200__A4 _00658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08011__B _02366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11971_ _00340_ clknet_leaf_39_wb_clk_i net47 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_99_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09686__A1 _02850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08489__A2 _02761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10296__A2 _04430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10922_ _04999_ _04700_ _05023_ _05024_ _04912_ _00355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XTAP_3978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_189_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10853_ _04708_ _04957_ _04958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_71_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10048__A2 _04173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_158_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08646__C1 as2650.stack\[11\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10784_ _02772_ _04891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_13_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_185_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_90_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11548__A2 _05556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11405_ _05455_ _05480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08413__A2 _02697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_181_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06424__A1 _00505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10220__A2 _00736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11336_ as2650.stack\[5\]\[7\] _05153_ _05154_ as2650.stack\[7\]\[7\] _05428_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_158_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_171_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10007__I _00749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11267_ _02613_ _05142_ _00759_ _05360_ _05361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_64_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08177__A1 _02325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10218_ _00789_ _04367_ _04368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09913__A2 _01619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11198_ _00439_ _05282_ _05285_ _05293_ _05294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__06727__A2 _00655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10149_ _00678_ _04301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_3_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07316__I _01751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06220__I _00677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09677__A1 _02055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11484__A1 _02028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_0 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_35_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11236__A1 as2650.stack\[1\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07360_ as2650.stack\[15\]\[8\] _01739_ _01795_ as2650.stack\[12\]\[8\] _01796_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_50_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11236__B2 as2650.stack\[3\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06311_ _00671_ _00762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_31_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07291_ _01726_ _01727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_176_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_30_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09030_ _03260_ _00227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_148_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_164_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06242_ _00698_ _00699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11701__CLK clknet_leaf_116_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_191_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06173_ _00631_ _00632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_172_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08404__A2 _02689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10211__A2 _00786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_1867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_176_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09932_ _04087_ _04088_ _04089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_67_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08168__A1 _02318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09863_ _03975_ _03976_ _04021_ _04022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07915__A1 _02181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08814_ _00955_ _00941_ _03061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09794_ _03951_ _03953_ _03954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07226__I _05724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06130__I _05771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08745_ _02394_ _02996_ _03003_ _03006_ _00196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05957_ _05789_ _05811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_38_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09668__B2 _03830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05941__A3 _05786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10278__A2 _02844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08676_ _01466_ _01433_ _02938_ _02947_ _02948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_54_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05888_ as2650.r0\[6\] _05742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_26_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08340__A1 _02525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07627_ net56 _02054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08891__A2 _03059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11227__A1 _02927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07558_ _00668_ _00855_ _01986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_50_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06509_ _00827_ _00950_ _00951_ _00952_ _00953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_195_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09840__A1 _02105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07489_ as2650.stack\[10\]\[12\] _01865_ _01872_ _01921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08643__A2 _02913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07896__I _02280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09228_ _03444_ _03446_ _03447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_158_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09159_ _03314_ _03378_ _03379_ _03380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_87_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_163_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06305__I _00755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10202__A2 _03697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06957__A2 _01396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_162_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11121_ _05216_ _05217_ _05218_ _05219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_174_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output70_I net70 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09616__I _03779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11052_ _05150_ _05151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_5111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_77_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_153_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10003_ _03917_ _04153_ _04154_ _04155_ _04158_ _04159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_7_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09659__A1 _00629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08676__B _02938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05932__A3 _05770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10269__A2 _04320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11466__A1 _00450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11954_ _00323_ clknet_leaf_19_wb_clk_i as2650.holding_reg\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_18_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07134__A2 _00666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10905_ _02212_ _04949_ _05008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10497__I _04608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11885_ _00254_ clknet_leaf_98_wb_clk_i as2650.stack\[4\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08882__A2 _03127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11218__A1 _05309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06893__A1 _01331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10836_ as2650.ivec\[3\] _04469_ _04941_ _04934_ _04642_ _04942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__11724__CLK clknet_leaf_113_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10767_ _02116_ _04789_ _04872_ _04874_ _00739_ _00350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_157_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09831__A1 _03987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06645__A1 _01086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06645__B2 _01088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10441__A2 _04076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10698_ _04801_ _04804_ _04805_ _04806_ _02824_ _04807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_157_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10729__B1 _04837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06948__A2 _01116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11319_ _03609_ _05189_ _05411_ _05412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_49_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08430__I _02709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11154__B1 _05249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06860_ _01008_ _01009_ _01301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_136_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06176__A3 _00633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08570__A1 _00630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06791_ _00423_ _01228_ _01232_ as2650.holding_reg\[2\] _01233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_114_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08530_ _01776_ _02798_ _02802_ _02803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_82_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11457__A1 _05517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09261__I _03470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08322__A1 _01934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08461_ _01026_ _02733_ _02734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_24_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07412_ _01821_ _01834_ _01843_ _01846_ _01847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA__11209__A1 _05216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06884__A1 as2650.holding_reg\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08392_ _02670_ _02682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07343_ _01743_ _01779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07274_ _01290_ _00848_ _01104_ _01710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__10432__A2 _02784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09013_ _03243_ _03067_ _03244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_192_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06225_ _00682_ _00683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_129_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08389__A1 _02678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_163_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06156_ _00614_ _00615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_172_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10196__A1 _04339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_1675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07061__A1 _01059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_1697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06087_ _00466_ _00545_ _00546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_82_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10803__C _00732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09915_ _00808_ _01693_ _04072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_144_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10499__A2 _05782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09846_ _03994_ _03998_ _04003_ _04004_ _04005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_63_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09777_ _02853_ _01302_ _03937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_132_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06989_ _01428_ _01429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_3027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11448__A1 _01223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08728_ _02412_ _02985_ _02991_ _02992_ _00193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_2304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08313__A1 _02609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08659_ net77 _02931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_14_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10120__A1 _04270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11206__I _01870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11670_ _00053_ clknet_leaf_130_wb_clk_i as2650.stack\[13\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10671__A2 _01738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10621_ as2650.stack\[1\]\[3\] _01815_ _01818_ as2650.stack\[0\]\[3\] as2650.stack\[2\]\[3\]
+ _01876_ _04732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XANTENNA__09813__A1 _03951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11897__CLK clknet_leaf_96_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_139_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10552_ _04658_ _04659_ _04663_ _04664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11620__A1 _04652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10423__A2 _04536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10266__B _03673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_194_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10483_ _04595_ _04596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_129_wb_clk_i clknet_4_0_0_wb_clk_i clknet_leaf_129_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_182_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07052__A1 _01420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05874__I _05727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11104_ _00774_ _05202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_123_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_172_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11035_ _05103_ _05134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08552__A1 _01598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11937_ _00306_ clknet_leaf_64_wb_clk_i net42 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10111__A1 _04256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08855__A2 _03101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07512__C1 _01942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11868_ _00237_ clknet_leaf_33_wb_clk_i as2650.r123_2\[2\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05913__I0 as2650.r123\[2\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10662__A2 _04748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09949__C _04105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10819_ _03740_ _04723_ _04925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_60_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09804__A1 _03933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11799_ _00182_ clknet_leaf_121_wb_clk_i as2650.stack\[15\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_140_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06618__A1 _01015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11611__A1 _04437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10414__A2 _04520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06094__A2 _00547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_173_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06010_ _00467_ _00468_ _00469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_31_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10178__A1 _02352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07043__A1 _05733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08791__A1 _02097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07594__A2 _02018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07961_ _02329_ _02279_ _02330_ _02281_ _00088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_87_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09700_ _02054_ _03790_ _03862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06912_ _01209_ _01211_ _01213_ _01220_ _01353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_68_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07892_ _01984_ _02270_ _02275_ _02282_ _00067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_68_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08543__A1 _02815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09631_ _03760_ _03794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_28_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06843_ _01150_ _01284_ _01285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_95_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09562_ _02039_ _03726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06774_ as2650.r123\[0\]\[2\] as2650.r123_2\[0\]\[2\] net51 _01216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_97_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_36_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08513_ as2650.stack\[5\]\[6\] _02785_ _01756_ as2650.stack\[4\]\[6\] _02786_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_110_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09493_ _03637_ _03643_ _03652_ _03659_ _03660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_97_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11026__I _05124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06857__A1 _01268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08444_ _02680_ _02717_ _02718_ _02719_ _00182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__10653__A2 _05767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08375_ _02198_ _02649_ _02254_ _02669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_149_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_162_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06609__A1 _01033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07326_ _01752_ _01762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__11602__A1 _02764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08335__I _02627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09271__A2 _03465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07282__A1 _05677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07257_ _01282_ _01690_ _01694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_136_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06208_ _00666_ _00667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_121_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05832__A2 _05685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07188_ _01536_ _01561_ _01625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_121_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10169__A1 _00546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09594__C _03757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_191_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07034__A1 _01316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07034__B2 _01319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06139_ _00597_ _00598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10533__C _04645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07585__A2 _02012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_48_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07337__A2 _01772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09829_ _02612_ _01474_ _03988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_100_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10341__A1 _00460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output33_I net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_161_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11722_ _00105_ clknet_leaf_4_wb_clk_i as2650.stack\[12\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_54_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_180_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11653_ _00036_ clknet_leaf_135_wb_clk_i as2650.stack\[13\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05869__I as2650.r0\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06863__A4 _00906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10604_ _03150_ _00896_ _04610_ _04714_ _04715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__10708__C _04109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout82 net83 net82 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout93 net30 net93 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_126_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11584_ _01462_ _02833_ _05628_ _04062_ _05629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_156_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10535_ _02057_ _02039_ _02070_ _04647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_13_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10466_ _03726_ _04533_ _04530_ _04579_ _04580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_142_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_clkbuf_leaf_29_wb_clk_i_I clknet_4_7_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10397_ _04481_ _04511_ _04512_ _04506_ _00342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
Xclkbuf_3_6_0_wb_clk_i clknet_0_wb_clk_i clknet_3_6_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_124_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08773__A1 _03020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11372__A3 _02664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11109__B1 _05204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10580__A1 as2650.stack\[14\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10580__B2 as2650.stack\[12\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_0_wb_clk_i_I wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_97_wb_clk_i clknet_4_9_0_wb_clk_i clknet_leaf_97_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_77_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08525__A1 _02789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11018_ _00963_ _04319_ _03745_ _00647_ _05117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_65_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11555__B _04225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_26_wb_clk_i clknet_4_5_0_wb_clk_i clknet_leaf_26_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_64_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_52_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06839__A1 _01252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10635__A2 _04701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06490_ _00933_ _00934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_59_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_166_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10685__I _01291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11721__D _00104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_68_wb_clk_i_I clknet_4_9_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08160_ as2650.stack\[7\]\[8\] _02488_ _02490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_158_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08155__I _02033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09253__A2 _03470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10399__A1 _02347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07111_ _05758_ _01217_ _01549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_147_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_119_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06067__A2 _00522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10938__A3 _04949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08091_ _02435_ _02436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07042_ _01432_ _00871_ _01481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07927__C _02306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07016__A1 _01138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08764__A1 _02415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_192_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06403__I _00667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08993_ _03033_ _03217_ _03227_ _03229_ _00221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_87_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10571__A1 as2650.stack\[5\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10571__B2 as2650.stack\[4\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07944_ _02277_ _02319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_9_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09714__I net89 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11465__B _05221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07875_ as2650.stack\[12\]\[14\] _02251_ _02267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_21_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06826_ _01266_ _01267_ _01268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09614_ _03777_ _03731_ _03778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__10874__A2 _03733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09545_ _02556_ _03708_ _03709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06757_ _01199_ _01200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08819__A2 _00995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_129_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09476_ _03639_ _03640_ _03642_ _03643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__10626__A2 _02782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_184_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06688_ _00541_ _00812_ _01130_ _01131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_51_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09492__A2 _03653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08493__C _02584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08427_ _02706_ _02707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_145_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08358_ _02516_ _02646_ _02652_ _02656_ _00159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_177_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_7_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07255__A1 _01601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06058__A2 _00516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07309_ _01744_ _01745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_138_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08289_ _02582_ _02337_ _02597_ _02598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_165_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10320_ _04450_ as2650.holding_reg\[6\] _04425_ _04451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_152_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07007__A1 _01442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10251_ _04395_ _04392_ _04396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_124_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07558__A2 _00855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08755__A1 _02405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07409__I _01775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06313__I _00656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10182_ _04332_ _04333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10562__A1 _00895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09624__I _02055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10314__A1 _04428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06469__B _00914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10865__A2 _04967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07730__A2 _02149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_102_wb_clk_i_I clknet_4_9_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_163_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08286__A3 _02573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11705_ _00088_ clknet_leaf_114_wb_clk_i as2650.stack\[10\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11290__A2 _01619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11636_ _00019_ clknet_leaf_39_wb_clk_i as2650.r123\[1\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_129_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_168_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07246__A1 _01341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06049__A2 _00507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11567_ _01327_ _02880_ _05613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07246__B2 _01498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11042__A2 _01032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08994__A1 as2650.stack\[7\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10518_ as2650.stack\[9\]\[1\] _01829_ _01826_ as2650.stack\[8\]\[1\] _04631_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_143_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08703__I _02705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11498_ as2650.r123\[3\]\[6\] _05551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_155_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06651__C _01094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10449_ _00879_ _00827_ _04563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_171_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07549__A2 _01910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10002__B1 _00818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11345__A3 _05436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06223__I _00562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_112_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10553__A1 _04652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_174_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05990_ _00448_ _05700_ _00449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06509__B1 _00951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05980__A1 _00437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09171__A1 _03388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07660_ _01905_ _02084_ _02085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__10856__A2 _04173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_38_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06611_ _00970_ _00987_ _00995_ _01055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_81_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07591_ _01987_ _02019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_34_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11808__CLK clknet_leaf_5_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07989__I _02356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09330_ _02632_ _03533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_94_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10608__A2 _05767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06542_ _00537_ _00631_ _00986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_34_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10629__B _04739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09261_ _03470_ _03478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__06288__A2 _00740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07485__A1 as2650.stack\[3\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06473_ _00512_ _00811_ _00791_ _00919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__11281__A2 _01934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08212_ _02527_ _02522_ _02523_ _02528_ _00141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_53_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09192_ _03395_ _03399_ _03412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_159_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09226__A2 _02223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08029__A3 _02388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08143_ as2650.stack\[8\]\[10\] _02477_ _02478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__11033__A2 _05131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08985__A1 _03020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08074_ _02418_ _02425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08985__B2 _03223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07025_ net1 _01464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_162_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10544__A1 _04654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06212__A2 _00670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_102_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08976_ _03204_ _03215_ _00218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_4806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_152_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07960__A2 _02278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_57_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_102_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07927_ _02304_ _02207_ _02308_ _02306_ _00076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_4839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_99_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10847__A2 _04947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07858_ _02255_ _02256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_60_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07712__A2 _01772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06809_ _01250_ _01251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_16_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07789_ _02200_ _02201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_38_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09528_ _02017_ _03692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09465__A2 _03627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_1892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06279__A2 _00732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09459_ _03561_ _03627_ _03628_ _03629_ _00287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XPHY_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08673__B1 _02836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11272__A2 _05302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__11214__I _01879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_16_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_164_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06308__I _00758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_177_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07228__A1 _01664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11421_ _03565_ _05487_ _05490_ _05491_ _00387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__11024__A2 _05118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_124_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_137_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_177_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11352_ _05413_ _05427_ _05434_ _05443_ _05148_ _05444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_158_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_193_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10274__B _04412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10783__A1 _04811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_192_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10303_ _02855_ _04437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_101_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_152_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06451__A2 _00896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11283_ _05373_ _05376_ _05377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08728__A1 _02412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10234_ _04374_ _00901_ _04375_ _04382_ _04383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_106_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08728__B2 _02992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10535__A1 _02057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10165_ _04313_ _04315_ _04316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05882__I _05712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09354__I _03545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07951__A2 _02319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10096_ net67 _01608_ _04249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_48_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09153__B2 _03163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09303__B _03493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10998_ _00799_ _05671_ _05097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07602__I _02029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11263__A2 _01518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_143_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_160_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07219__A1 _01631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11015__A2 _05113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11619_ _02050_ _05657_ _05659_ _00712_ _00417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_121_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08967__A1 _01700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_190_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08433__I _02705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10774__A1 _02125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06442__A2 _00883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08719__A1 as2650.stack\[15\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_41_wb_clk_i clknet_4_6_0_wb_clk_i clknet_leaf_41_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10526__A1 _04622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08830_ _01026_ _03076_ _03077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07493__B _01924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08761_ _02412_ _03011_ _03016_ _03017_ _00201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_57_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05973_ _05792_ _00432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09144__A1 _05742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07712_ _02131_ _01772_ _02132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10829__A2 _04934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08692_ _00865_ _02807_ _02964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_26_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07643_ net89 _02069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_38_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07574_ _01819_ _02002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_78_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_81_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09313_ _02388_ _02438_ _03218_ _03520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_94_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06525_ _00944_ _00954_ _00968_ _00969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_22_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11254__A2 _05348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07458__B2 as2650.stack\[5\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09244_ _03446_ _03462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06456_ _00720_ _00725_ as2650.cycle\[12\] as2650.cycle\[7\] _00902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_107_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09175_ _05758_ _02233_ _03396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11006__A2 _00648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06387_ _00825_ _00832_ _00833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_108_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08126_ as2650.stack\[0\]\[7\] _02445_ _02435_ _02464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__10806__C _04912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08057_ _02409_ _02406_ _02410_ _02411_ _00103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xoutput15 net84 io_oeb[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_162_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput26 net26 io_out[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput37 net37 io_out[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_07008_ _01251_ _01429_ _01447_ _01293_ _01448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_122_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput48 net48 la_data_out[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput59 net86 la_data_out[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__10517__A1 _02780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_5315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11190__A1 _01028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07933__A2 _02227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_5359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08959_ _01596_ _03122_ _03125_ _03199_ _03200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_130_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09135__A1 _05750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_56_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11970_ _00339_ clknet_leaf_39_wb_clk_i net46 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_4669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09686__A2 _03803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10921_ as2650.ivec\[6\] _04972_ _04941_ _05002_ _04643_ _05024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XTAP_3968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07850__C _02047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10852_ _04946_ _04957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__07422__I _01795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10783_ _04811_ _04877_ _04890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_12_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08646__B1 _02795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08646__C2 _02799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_184_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07578__B _00956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05877__I as2650.r0\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09349__I _02644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11404_ as2650.stack\[9\]\[1\] _05478_ _05479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_172_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11335_ _05796_ _05282_ _05416_ _05426_ _05427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__06424__A2 _00834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07621__A1 _01984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11266_ _02837_ _02960_ _05359_ _02810_ _05360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_107_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10508__A1 _00929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_190_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08177__A2 _02500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09374__A1 _03565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10217_ net91 _02808_ _00496_ _00787_ _04367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_140_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11197_ _02842_ _03815_ _05291_ _05292_ _05293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_45_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07385__B1 _01819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07924__A2 _02197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10148_ _02225_ _04069_ _04299_ _04300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_95_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05935__A1 _05787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10079_ _04228_ _04232_ _04233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__12009__CLK clknet_leaf_117_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09677__A2 _01141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09812__I _02893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07688__A1 _02104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08885__B1 _03130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06360__A1 _00543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_1 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__10179__B _03646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07332__I net70 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11236__A2 _05162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06310_ _00757_ _00696_ _00588_ _00760_ _00761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_31_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07290_ _01290_ _01725_ _01104_ _01726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_148_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10995__A1 _01974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06241_ _00576_ _00698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10693__I _00444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07860__A1 _02197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_191_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06172_ _00536_ as2650.cycle\[1\] _00631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_117_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08163__I _02492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09601__A2 _01019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10747__A1 _04023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_1857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_1879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09931_ net36 net35 _03996_ _04088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_137_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07935__C _02158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08168__A2 _02489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09365__A1 _03558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09862_ _04006_ _04020_ _03883_ _04021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07915__A2 _02297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08813_ _00953_ _03055_ _03057_ _03059_ _03060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_98_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09793_ _03952_ _03902_ _03953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_189_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05956_ _05790_ _05757_ _05809_ _05769_ _05810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_113_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08744_ as2650.stack\[1\]\[1\] _03004_ _03005_ _03006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_27_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09668__A2 _03815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08675_ _02944_ _02945_ _02946_ _02947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_54_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05887_ _05735_ _05740_ _05741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_76_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07626_ _02052_ _02053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_14_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07557_ _01773_ _01985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_179_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06508_ _00489_ _00952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10435__B1 _04542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06103__A1 _00531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07488_ as2650.stack\[9\]\[12\] _01869_ _01758_ as2650.stack\[8\]\[12\] as2650.stack\[11\]\[12\]
+ _01740_ _01920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_50_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09840__A2 _01464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10986__A1 _00805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09227_ _03418_ _03422_ _03445_ _03446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06654__A2 _01097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06439_ _00884_ _00885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07398__B _01788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_148_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09158_ _03348_ _03371_ _03379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_87_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08109_ as2650.stack\[0\]\[3\] _02440_ _02451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06406__A2 _00657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09089_ _01643_ _03309_ _03311_ _03312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__10202__A3 _04346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11120_ as2650.stack\[2\]\[1\] _05212_ _05157_ as2650.stack\[0\]\[1\] _05218_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_89_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09356__A1 as2650.stack\[3\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11051_ _01992_ _05149_ _05150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_5101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_104_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_output63_I net63 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08022__B _02356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11163__A1 as2650.stack\[2\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10002_ _04157_ _03872_ _00818_ _04131_ _03925_ _04158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_118_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_191_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_190_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10910__A1 _04609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09659__A2 _03821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09632__I net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08676__C _02947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11953_ _00322_ clknet_leaf_20_wb_clk_i as2650.holding_reg\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10269__A3 _04407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11466__A2 _02768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08331__A2 _02636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_189_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10904_ _05001_ _05007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_3798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11884_ _00253_ clknet_leaf_103_wb_clk_i as2650.stack\[4\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06893__A2 _01333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08619__B1 _02871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10835_ _02557_ _04941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_25_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06991__I _01297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_185_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10766_ as2650.ivec\[1\] _04470_ _04841_ _04845_ _04873_ _04874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_125_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07842__A1 _02239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10697_ _00444_ _04806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_145_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11318_ _00824_ _05394_ _05401_ _05410_ _05278_ _05411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_141_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10462__B _03738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11249_ _05340_ _05343_ _05344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_171_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11154__A1 _03138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_95_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08945__I1 _01458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06231__I _00688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10901__A1 _03820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06790_ _00421_ _01064_ _01231_ _00828_ _01232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_95_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06581__A1 _00745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11457__A2 _03484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08322__A2 _01769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10665__B1 _01756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08460_ _02732_ _02727_ _02733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_63_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07530__B1 _01944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07411_ _01845_ _01846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_63_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08391_ _02666_ _02681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_162_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06884__A2 _00829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07997__I _02059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07342_ _01763_ _01767_ _01777_ _01778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_108_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_176_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07273_ as2650.r123\[0\]\[0\] _01709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_104_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07833__A1 _02222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11699__CLK clknet_leaf_123_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_148_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09012_ _05696_ _00826_ _03243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08107__B _02446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06224_ _00638_ _00681_ _00682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_164_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08389__A2 _02667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_1643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06155_ _00492_ _00503_ _05701_ _00614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA_clkbuf_4_1_0_wb_clk_i_I clknet_3_0_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10196__A2 _04345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11393__A1 _02684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08621__I _02893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06086_ _00543_ _00544_ _00545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_105_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09338__A1 _03239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09914_ _04026_ _04029_ _04070_ _04071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_132_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11145__A1 _02814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08010__A1 as2650.stack\[14\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09845_ _03776_ _04004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09776_ _03933_ _03935_ _03936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_3006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06988_ _01299_ _01424_ _01425_ _01426_ _01427_ _01428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XTAP_3017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_160_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08727_ _02461_ _02712_ _02969_ _02992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_2305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11448__A2 _03454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05939_ _05757_ _05792_ _05763_ _05769_ _05793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_96_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_160_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09510__A1 _00622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08068__I _02419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08658_ net85 _02930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_1615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_4_8_0_wb_clk_i clknet_3_4_0_wb_clk_i clknet_4_8_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_1626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07609_ net90 _02037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_41_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08589_ _02860_ _02613_ _02861_ _02862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_54_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10620_ _01734_ _04729_ _04730_ _04731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__10959__A1 _02229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10547__B _04588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09813__A2 _03837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07700__I _05687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10551_ _04590_ _04661_ _04662_ _02334_ _04663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_122_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11620__A2 _04399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10266__C _04405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10482_ _00443_ _04595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09577__A1 _00638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_19_wb_clk_i_I clknet_4_5_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09627__I net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11103_ _04275_ _01127_ _05201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11809__D _00192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09329__A1 _03037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11136__A1 _05221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06051__I _05676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11034_ _02028_ _02589_ _02724_ _05133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08001__A1 _02051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06938__I0 as2650.r123\[0\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08687__B _02958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08552__A2 _02590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06563__A1 _01001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09362__I _02076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11439__A2 _03374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_185_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11936_ _00305_ clknet_leaf_61_wb_clk_i net41 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07512__B1 _01941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07512__C2 as2650.stack\[1\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11867_ _00236_ clknet_leaf_33_wb_clk_i as2650.r123_2\[2\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11841__CLK clknet_leaf_102_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10818_ _04709_ _04921_ _04923_ _02334_ _04924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__08706__I _02059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09804__A2 _03963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07610__I _02037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11798_ _00181_ clknet_leaf_120_wb_clk_i as2650.stack\[15\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_41_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10749_ _00445_ _04846_ _04856_ _02901_ _04857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__11611__A2 _05575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10414__A3 _04523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11991__CLK clknet_leaf_26_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06094__A3 _00552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_173_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_145_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_192_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10178__A2 _00899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07043__A2 _00962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08240__A1 _00650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_142_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08791__A2 _03029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07960_ as2650.stack\[10\]\[14\] _02278_ _02330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_142_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06911_ _01202_ _01221_ _01352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07891_ _02276_ _02279_ _02281_ _02282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_151_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09740__A1 _03893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09630_ _00538_ _03793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08543__A2 _01032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06842_ _01282_ _01157_ _01284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06554__A1 _00921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06773_ _01209_ _01211_ _01214_ _01215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09561_ _03724_ _03725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_23_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_97_wb_clk_i_I clknet_4_9_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08512_ _02784_ _02785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_77_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09492_ _02568_ _03653_ _03656_ _03658_ _03659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_36_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06857__A2 _01255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08443_ as2650.stack\[15\]\[12\] _02714_ _02719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08374_ as2650.stack\[2\]\[8\] _02666_ _02668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08059__A1 as2650.stack\[12\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09256__B1 _03473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08616__I _01711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07325_ _01757_ _01761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07806__A1 _02189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11602__A2 _02740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07256_ _01692_ _01693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_137_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06207_ _00665_ _00666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07187_ _01536_ _01561_ _01624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_117_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10169__A2 _02599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09447__I _02534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06138_ _00594_ _00596_ _00597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07034__A2 _01453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11198__B _05285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08231__A1 as2650.stack\[5\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_156_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07585__A3 _00576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06069_ net5 _00528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__06793__A1 as2650.holding_reg\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09731__A1 _03887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09828_ _03943_ _03985_ _03944_ _03986_ _03987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_86_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10341__A2 _04457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09759_ _03908_ _03919_ _03920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_100_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output26_I net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09910__I _03719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11721_ _00104_ clknet_leaf_5_wb_clk_i as2650.stack\[12\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_154_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11652_ _00035_ clknet_leaf_2_wb_clk_i as2650.stack\[13\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10603_ _04391_ _04587_ _04714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xfanout83 net84 net83 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_128_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11583_ _05356_ _05627_ _05241_ _05628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xfanout94 net53 net94 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_122_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10534_ _03876_ _02055_ _02038_ _04646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_10_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08470__A1 _00763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10465_ _03916_ _04578_ _04579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_124_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08222__A1 as2650.stack\[5\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08261__I _00602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10396_ net22 _04487_ _04512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_123_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09970__A1 _03849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08773__A2 _03022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11109__A1 _04460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11109__B2 _03782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10580__A2 _04681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_131_wb_clk_i_I clknet_4_0_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09722__A1 _02071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11017_ _05100_ _05107_ _05115_ _05116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__09306__B _03493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06536__A1 as2650.addr_buff\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11127__I _01811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10031__I _04173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08289__A1 _02582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_66_wb_clk_i clknet_4_12_0_wb_clk_i clknet_leaf_66_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_3381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10096__A1 net67 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06839__A2 _01157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11919_ _00288_ clknet_leaf_96_wb_clk_i as2650.stack\[5\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08436__I _02705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07340__I _01775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09789__A1 _02859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07110_ _05750_ _01379_ _01548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_53_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08090_ _02422_ _02435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_174_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07264__A2 _01700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06067__A3 _00525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08461__A1 _01026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07041_ _01432_ _00830_ _01479_ _01480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_122_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_173_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11348__A1 _05209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10634__C _04744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07016__A2 _05793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08213__A1 _02030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11737__CLK clknet_leaf_108_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09961__A1 _00792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08764__A2 _03011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08992_ as2650.stack\[7\]\[2\] _03228_ _03225_ _03229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_173_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10571__A2 _02913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07943_ _02206_ _02318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_155_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09713__A1 _00523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_68_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07874_ _02231_ _02263_ _02264_ _02266_ _00065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_56_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11520__A1 _05556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11520__B2 _03780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09613_ _03776_ _03777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06825_ _05745_ _05767_ _05768_ _05739_ _01267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_99_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09544_ _05703_ _00458_ _00949_ _03672_ _03708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_06756_ _01198_ _01199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_70_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_93_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08819__A3 _03054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10087__A1 net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06687_ _00993_ _01130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09475_ _03641_ _03642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_149_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08426_ _02705_ _02706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08357_ as2650.stack\[3\]\[10\] _02655_ _02656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_138_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11587__A1 _02101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07308_ _01743_ _01744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07255__A2 _01011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08452__A1 _02723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08288_ _05696_ _02335_ _02596_ _02597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_20_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06463__B1 _00901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07239_ _01674_ _01675_ _01676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_118_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11339__A1 as2650.stack\[0\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10250_ as2650.addr_buff\[4\] _04395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06215__B1 _00673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08755__A2 _03011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10181_ _04331_ _04332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_160_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06766__A1 _00999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10560__B _04671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06518__A1 _00478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10314__A2 _04397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11511__A1 _05150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07425__I _01791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07191__A1 _01539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_28_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12042__CLK clknet_opt_1_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09640__I _03766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11391__B _05468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11704_ _00087_ clknet_leaf_114_wb_clk_i as2650.stack\[10\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08691__A1 _02811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07160__I _01597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11635_ _00018_ clknet_leaf_27_wb_clk_i as2650.r123\[1\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11578__A1 _01983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11566_ _01576_ _01583_ _02875_ _01679_ _05612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_11_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10517_ _02780_ _04625_ _04629_ _04630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_11497_ _05550_ _00404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_155_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_113_wb_clk_i clknet_4_2_0_wb_clk_i clknet_leaf_113_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_155_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06504__I _00487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10448_ _02038_ _04560_ _05703_ _04562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_170_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10002__A1 _04157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10026__I net39 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10002__B2 _04131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09943__A1 _04087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08746__A2 _02998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10379_ _04489_ _04497_ _04498_ _00338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_112_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09815__I _00727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_152_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12049_ _00418_ clknet_leaf_18_wb_clk_i net29 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_61_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11285__C _05185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06509__A1 _00827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10856__A3 _04930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08875__B _03072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06610_ _01013_ _01023_ _01053_ _01054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_25_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07590_ _02004_ _02015_ _02017_ _02018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_94_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06541_ as2650.cycle\[9\] _00985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__10696__I _04792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09260_ _03459_ _03472_ _03476_ _03477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06472_ _00900_ _00909_ _00917_ _00918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_107_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08682__A1 _02597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07485__A2 _01862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08211_ as2650.stack\[6\]\[14\] _02507_ _02528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09191_ _03382_ _03403_ _03411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_163_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09226__A3 _03423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08029__A4 _02023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08142_ _02466_ _02477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10645__B _04754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10241__A1 _04186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08073_ _02314_ _02420_ _02421_ _02424_ _00106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_11_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_161_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07024_ _01433_ _05803_ _01463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_162_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_134_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09934__A1 _00719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_192_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06748__A1 _01060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09725__I net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_5508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08975_ _01658_ _03177_ _03214_ _03099_ _03215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_9_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_64_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_102_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07926_ as2650.stack\[11\]\[9\] _02307_ _02308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_4829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_116_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09162__A2 _03366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_84_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07857_ _02154_ _02136_ _02254_ _02255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_56_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06808_ _00970_ _00987_ _00995_ _01250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_28_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06920__A1 _01357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07788_ _02199_ _02200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_71_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09527_ _00577_ _00579_ _00581_ _00567_ _03691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_06739_ _01180_ _01181_ _01182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_129_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08673__A1 _02848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09458_ as2650.stack\[5\]\[4\] _03620_ _03621_ _03629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08673__B2 _02940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11902__CLK clknet_leaf_73_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__10480__A1 _00780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08409_ _02688_ _02695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09389_ _02045_ _03579_ _02523_ _03580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_138_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11420_ _02110_ _05462_ _05472_ _05491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_142_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08425__A1 _02154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11024__A3 _05122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07848__C _02047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10232__A1 _03877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08976__A2 _03215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11351_ _05221_ _05442_ _05443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06987__A1 _01309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_152_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10783__A2 _04877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10302_ _04426_ _04435_ _04436_ _00323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_180_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06324__I _00774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11282_ _05298_ _05374_ _05375_ _05376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_152_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09925__A1 _01610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08728__A2 _02985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10233_ _03655_ _04378_ _04380_ _04381_ _04382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_161_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06739__A1 _01180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10535__A2 _02039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10164_ _00938_ _02333_ _04314_ _04315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_117_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10095_ _00719_ _04245_ _04247_ _03995_ _03777_ _04248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_0_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05962__A2 _05754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10299__A1 _02618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09153__A2 _03342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06994__I net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06911__A1 _01202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11405__I _05455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10997_ _05077_ _04701_ _05096_ _05076_ _00358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_90_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_182_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09861__B1 _03916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08416__A1 _02678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11618_ _05413_ _04638_ _05657_ _05658_ _05659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_89_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10223__A1 _00565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11549_ _05588_ _05595_ _04501_ _05596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_171_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06978__A1 _01094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10184__C _04334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06442__A3 _00660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09916__A1 _04071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08719__A2 _02972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_4_6_0_wb_clk_i_I clknet_3_3_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_124_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10526__A2 _04638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_98_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_4_10_0_wb_clk_i clknet_3_5_0_wb_clk_i clknet_4_10_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_98_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08760_ _02461_ _02695_ _02995_ _03017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05972_ _05771_ _05773_ _00430_ _00431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XTAP_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05953__A2 _05806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_81_wb_clk_i clknet_4_8_0_wb_clk_i clknet_leaf_81_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_66_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07711_ net59 _02131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08691_ _02811_ _02962_ _02963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_66_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08498__A4 _02770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07642_ as2650.stack\[13\]\[2\] _02025_ _02068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_54_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06902__A1 _01342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11925__CLK clknet_leaf_62_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06753__I1 _01195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11239__B1 _05163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07573_ _02000_ _02001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09312_ _03518_ _03519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06524_ _00955_ _00957_ _00967_ _00968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_22_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07458__A2 _01858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09852__B1 _03997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09243_ _03439_ _03443_ _03461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__10462__A1 _03749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06455_ _00862_ _00557_ _00901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_72_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09174_ _03323_ _03394_ _03361_ _03362_ _03395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_147_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06386_ _00826_ _00827_ _00767_ _00831_ _00832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_21_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11006__A3 _00870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08125_ _02381_ _02442_ _02463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_162_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08056_ _02177_ _02258_ _02385_ _02411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_116_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput16 net16 io_oeb[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput27 net27 io_out[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_190_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07007_ _01442_ _01446_ _01288_ _01447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_137_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09907__A1 _04023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput38 net38 io_out[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__09907__B2 _03977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput49 net49 la_data_out[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_89_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08958_ _03197_ _03198_ _03122_ _03199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_88_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_102_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05944__A2 _05793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07909_ _02091_ _02292_ _02294_ _02295_ _00071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_44_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08889_ _03059_ _03134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_3925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_99_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_99_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10920_ _03662_ _05002_ _05021_ _05022_ _03832_ _05023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XTAP_3958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08894__A1 _03138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_29_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10851_ _04167_ _04228_ _04955_ _04956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_38_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08646__A1 as2650.stack\[9\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10782_ _02952_ _04097_ _04888_ _04889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_25_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08646__B2 as2650.stack\[8\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_188_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__10453__A1 _00520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_164_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08534__I _02806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10285__B _00966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10205__A1 _00580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08949__A2 _03190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11403_ _05475_ _05478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_184_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_177_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11402__B1 _05474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09071__A1 _03214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10756__A2 _04863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11334_ _05424_ _05425_ _05426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06054__I _00492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07621__A2 _01998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06989__I _01428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11265_ _02812_ _05358_ _05359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_180_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10508__A2 _02727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10216_ _04314_ _04365_ _03755_ _04366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_106_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09374__A2 _03562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11196_ _01269_ _02866_ _03653_ _02856_ _05292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__07385__A1 as2650.stack\[5\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07385__B2 as2650.stack\[4\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10147_ _04287_ _04297_ _04298_ _04299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_62_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11948__CLK clknet_4_14_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10078_ _04217_ _04231_ _04232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_47_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08885__A1 _01206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07688__A2 _02110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08709__I _02710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08885__B2 as2650.r123_2\[1\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06735__I1 _00434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10692__A1 _02105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06360__A2 _00806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__10179__C _03781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06229__I _00562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09968__C _04082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_188_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10444__A1 _04376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06240_ _00696_ _00697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_15_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07860__A2 _02252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05871__A1 _05688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06171_ _00629_ _00630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_106_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09062__A1 _03189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_156_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09930_ net37 _04087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_131_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09861_ _04007_ _03724_ _03916_ _04019_ _04020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_113_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08812_ _03058_ _03059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_112_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10214__I _04363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09792_ net33 _03952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08743_ _02693_ _03005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05955_ _05784_ _05809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_100_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07128__A1 as2650.holding_reg\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08674_ _00626_ _01601_ _01138_ _01042_ _01460_ _01435_ _02946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_05886_ _05719_ _05737_ _05738_ _05739_ _05740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_26_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07523__I _01459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10683__A1 _04007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07625_ _02035_ _02052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06139__I _00597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07556_ _01983_ _01984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_41_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10435__A1 as2650.stack\[15\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10884__I _04987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06507_ _00650_ _00951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_22_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10435__B2 as2650.stack\[14\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_194_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06103__A2 _00561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07487_ _01917_ _01918_ _01846_ _01919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_42_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05978__I _05769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09226_ _01663_ _02223_ _03423_ _03445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_107_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06438_ _00663_ _00884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09428__I0 as2650.ivec\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05862__A1 _05708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09157_ _03348_ _03371_ _03378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_166_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09053__A1 _01926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09894__B _04051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06369_ _00607_ _00559_ _00815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_159_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08108_ _02399_ _02436_ _02448_ _02450_ _00115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_09088_ _01550_ _03310_ _03311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_120_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08800__A1 _02461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10202__A4 _04351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_150_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08039_ as2650.stack\[12\]\[1\] _02396_ _02397_ _02398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_194_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06602__I _01035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11050_ _02131_ _01990_ _05149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_118_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11163__A2 _05212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10001_ _04156_ _04157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_131_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output56_I net56 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_184_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_4445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11952_ _00321_ clknet_4_5_0_wb_clk_i as2650.holding_reg\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_123_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10903_ _04709_ _05004_ _05005_ _04419_ _05006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_3788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11883_ _00252_ clknet_leaf_103_wb_clk_i as2650.stack\[4\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_83_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08619__A1 _02778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10834_ _04161_ _04934_ _04939_ _03780_ _04940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA_clkbuf_leaf_48_wb_clk_i_I clknet_4_13_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08619__B2 _02891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09292__A1 as2650.stack\[2\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10765_ _04642_ _04873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__05888__I as2650.r0\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07842__A2 _02214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09419__I0 as2650.ivec\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10696_ _04792_ _04805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_31_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_185_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10729__A2 _04793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11317_ _05185_ _05409_ _05410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_173_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09309__B _03493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07608__I _02035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11770__CLK clknet_leaf_92_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11248_ _05160_ _05341_ _05342_ _05343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_136_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11154__A2 _02815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11179_ _05265_ _05275_ _05276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_132_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10901__A2 _04262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06581__A2 _01024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_149_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10665__A1 as2650.stack\[7\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10665__B2 as2650.stack\[4\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07530__B2 as2650.stack\[6\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07410_ _01844_ _01845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_23_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08390_ _02226_ _02680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_36_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09698__C _03859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07341_ _01776_ _01777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07499__B _01930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08086__A2 _02427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09283__A1 _03000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10968__A2 _05063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11090__A1 _03974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08174__I _02488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07272_ _01659_ _01708_ _00021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07833__A2 _02237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05844__A1 _05697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09011_ _03050_ _03233_ _03241_ _03242_ _00226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_178_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06223_ _00562_ _00681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09035__A1 _03129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_191_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06154_ _00612_ _00613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_1655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11393__A2 _05467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06085_ as2650.cycle\[13\] _00535_ _00544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_171_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08123__B _02435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09913_ _01610_ _01619_ _04070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09338__A2 _02634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11145__A2 _00842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09844_ _04000_ _04002_ _04003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_113_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08010__A2 _02362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09733__I _03762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_189_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09775_ _03906_ _03934_ _03935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_74_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06987_ _01309_ _01259_ _01427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_3007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08726_ as2650.stack\[15\]\[6\] _02978_ _02991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05938_ _05784_ _05792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10656__A1 _04763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09510__A2 _00911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08657_ _01772_ _01043_ _01142_ _01771_ _02929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_15_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05869_ as2650.r0\[7\] _05723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_81_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07608_ _02035_ _02036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_42_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08588_ _02826_ _02861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10408__A1 _00602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_180_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07539_ as2650.stack\[11\]\[14\] _01959_ _01735_ _01969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_167_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11643__CLK clknet_leaf_32_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06088__A1 _00541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10959__A2 _00628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10550_ _00780_ _04648_ _04662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_139_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09209_ _03426_ _03428_ _03429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__05835__A1 _05687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09026__A1 _00838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_167_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10481_ _04590_ _04592_ _04593_ _02334_ _04594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_87_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09577__A2 _00893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08812__I _03058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11793__CLK clknet_leaf_86_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07588__A1 _00568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07428__I _01739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08033__B _02264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11102_ _00774_ _05200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_150_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06332__I _00458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_121_wb_clk_i_I clknet_4_0_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_85_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11033_ net78 _05131_ _05132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_150_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07872__B _02264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08001__A2 _02357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10344__B1 _04458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06938__I1 as2650.r123_2\[0\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06012__A1 _00466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10895__A1 _04223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06563__A2 _00966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11825__D _00208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07760__A1 _02091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08259__I _02567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_4_wb_clk_i_I clknet_4_1_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10647__A1 _04709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11935_ _00304_ clknet_leaf_64_wb_clk_i net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_27_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07512__A1 as2650.stack\[3\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11866_ _00235_ clknet_leaf_34_wb_clk_i as2650.r123_2\[2\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_150_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10817_ _04808_ _04922_ _04923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_53_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09265__A1 _03439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11797_ _00180_ clknet_leaf_120_wb_clk_i as2650.stack\[15\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_9_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10748_ _04802_ _04855_ _04856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06507__I _00650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10414__A4 _04527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10679_ _02094_ _04701_ _04788_ _04645_ _00348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_173_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09818__I _00748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07579__A1 _00513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08240__A2 _02546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06242__I _00698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06251__A1 _00482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06251__B2 _00707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08528__B1 _02795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06910_ _01324_ _01350_ _01000_ _01351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_96_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07890_ _02280_ _02281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_110_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06003__A1 _00460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10920__C _03832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06841_ _01255_ _01256_ _01282_ _01283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XANTENNA__09740__A2 _03900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08543__A3 _01454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10886__A1 _04725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06554__A2 _00997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07751__A1 _02067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09560_ _00748_ _02866_ _03724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_110_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06772_ _01213_ _01214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_83_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08511_ _01749_ _02784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_184_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09491_ _03657_ _02546_ _03658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_58_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11666__CLK clknet_leaf_121_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08442_ _02710_ _02718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_169_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09502__B _00648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07801__I net66 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08373_ _02666_ _02667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09256__B2 _03177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10367__C _04405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07324_ _01735_ _01748_ _01759_ _01760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_143_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06417__I _00862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07806__A2 _02214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11602__A3 _03638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07255_ _01601_ _01011_ _01688_ _01426_ _01691_ _01692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__09008__A1 _03047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07282__A3 _01717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06206_ _00664_ _00665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_121_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07186_ _01564_ _01623_ _00020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10383__B _04501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10169__A3 _04319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06137_ _00595_ _00587_ _00596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_172_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08231__A2 _02538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10574__B1 _02914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_160_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06068_ _00475_ _00499_ _00509_ _00526_ _00527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XANTENNA__06793__A2 _00655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07990__A1 _02151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05991__I _00449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09827_ _03978_ _01444_ _03986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10877__A1 _04808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_59_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09731__A2 _03891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09758_ _03838_ _03864_ _03918_ _03919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_21_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08709_ _02710_ _02979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09689_ _03797_ _01159_ _01160_ _03798_ _03799_ _03851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_4
XTAP_2136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11720_ _00103_ clknet_leaf_5_wb_clk_i as2650.stack\[12\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07711__I net59 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output19_I net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_145_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11651_ _00034_ clknet_leaf_134_wb_clk_i as2650.stack\[13\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_147_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10277__C _04405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07258__B1 _01688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10602_ _04709_ _04711_ _04712_ _04419_ _04713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_126_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11582_ _05138_ _04446_ _05626_ _05627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
Xfanout84 net15 net84 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_183_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_167_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10533_ _02057_ _04531_ _04644_ _04645_ _00345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__10801__A1 _02621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08470__A2 _02742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08542__I _02814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06481__A1 as2650.cycle\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10464_ _03726_ _04535_ _02758_ _04553_ _04577_ _04578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_142_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_170_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10395_ _03609_ _04483_ _04510_ _04511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_123_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08222__A2 _02536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06233__A1 _00553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06062__I _00520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07430__B1 _01863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07430__C2 as2650.stack\[1\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11109__A2 _03679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11016_ _00880_ _05109_ _05114_ _05115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__10868__A1 as2650.ivec\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09722__A2 _03725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10868__B2 _04947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06536__A2 _00979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_187_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_185_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09486__A1 _00502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08289__A2 _02337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11918_ _00287_ clknet_leaf_72_wb_clk_i as2650.stack\[5\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11293__A1 net85 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06839__A3 _01253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_178_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09238__A1 _03189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11849_ _00009_ clknet_4_12_0_wb_clk_i as2650.cycle\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_61_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11045__A1 _02845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06237__I as2650.cycle\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_leaf_35_wb_clk_i clknet_4_6_0_wb_clk_i clknet_leaf_35_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_105_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11596__A2 _05637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06681__B _01123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07040_ _01478_ _00830_ _01479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_146_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_127_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11348__A2 _05438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09410__A1 _02119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06224__A1 _00638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09961__A2 _01692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08991_ _03219_ _03228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_138_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07942_ _02314_ _02315_ _02316_ _02317_ _00082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_44_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09713__A2 _03827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10859__A1 _04794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07873_ as2650.stack\[12\]\[13\] _02260_ _02266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_29_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09612_ _00632_ _03776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_28_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06824_ _01265_ _01065_ _01266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_95_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09543_ _00747_ _00546_ _03645_ _03707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_55_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06755_ as2650.r123\[0\]\[1\] as2650.r123_2\[0\]\[1\] _05710_ _01198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_97_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09477__A1 _00928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07488__B1 _01758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09474_ _02823_ _03641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06686_ _00904_ _00965_ _01128_ _01129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_110_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07488__C2 _01740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10378__B _04301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07531__I _01900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_93_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08425_ _02154_ _02031_ _02664_ _02705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_24_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08356_ _02644_ _02655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_51_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06147__I _00605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07307_ _01741_ _01742_ _01743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__11587__A2 _05624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08287_ _00837_ _00481_ _02596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_192_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08452__A2 _00870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05986__I _00444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06463__A1 _00509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07238_ _01670_ _01675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06463__B2 _00908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_30_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_152_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11339__A2 _05210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07169_ net2 _01607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09401__A1 _03558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06215__A1 _00464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06215__B2 _00525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_191_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10180_ _00578_ _04331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_65_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06766__A2 _01196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11831__CLK clknet_leaf_27_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09407__B _03574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06518__A2 _00961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_189_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09921__I _04077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09468__A1 _03571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_182_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11275__A1 _05298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08537__I _02764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10617__A4 _04727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07441__I _01779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11703_ _00086_ clknet_leaf_115_wb_clk_i as2650.stack\[10\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_15_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11027__A1 _03794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11634_ _00017_ clknet_leaf_37_wb_clk_i as2650.r123\[1\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_42_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09796__C _02890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11578__A2 _05611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11565_ _02965_ _05521_ _05610_ _05611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_10_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05896__I as2650.r0\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06454__A1 _00468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10516_ _04626_ _04627_ _04628_ _04629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__08272__I _02580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06454__B2 _00899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11496_ as2650.r123\[3\]\[5\] _05550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_156_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10447_ _02038_ _04560_ _00441_ _04561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_67_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10002__A2 _03872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10378_ net45 _04494_ _04301_ _04498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_123_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09317__B _02640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12048_ _00417_ clknet_leaf_9_wb_clk_i net79 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_26_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06509__A2 _00950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07706__A1 _02126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07182__A2 _01619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09459__A1 _03561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10977__I _02235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06540_ _00970_ _00981_ _00983_ _00984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__11266__A1 _02837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08667__C1 _02076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_179_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07351__I _01786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06471_ _00910_ _00916_ _00917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_61_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08891__B _03113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08210_ _02236_ _02527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_60_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11018__A1 _00963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_194_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09190_ _03408_ _03409_ _03410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_37_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11704__CLK clknet_leaf_114_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08141_ _02318_ _02468_ _02474_ _02476_ _00122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_53_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08434__A2 _02712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11601__I _05608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_174_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06445__A1 _00557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10241__A2 _04388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08182__I _02196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08072_ _02423_ _02424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_179_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07023_ _01461_ _01462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__11854__CLK clknet_leaf_54_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08198__A1 _02516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09934__A2 _04086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07945__A1 as2650.stack\[10\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08974_ _01686_ _03178_ _03213_ _03214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_142_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_116_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07925_ _02155_ _02307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_57_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09698__A1 _03774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07856_ _01988_ _02254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_56_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06807_ _01094_ _01230_ _01241_ _01248_ _01249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_4
XFILLER_186_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07787_ _02198_ _01989_ _01995_ _02199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__06920__A2 _05775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11257__A1 _00775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09526_ _03688_ _03689_ _03690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06738_ _01173_ _01174_ _01178_ _01181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_43_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_169_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_149_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09457_ _03509_ _03617_ _03628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06669_ _01102_ _01107_ _01112_ _01113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XPHY_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09897__B _04051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08673__A2 _01234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11009__A1 _02349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08408_ _02663_ _02690_ _02691_ _02694_ _00171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_12_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10480__A2 _04581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09388_ _02506_ _03579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_71_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08339_ as2650.stack\[4\]\[13\] _02636_ _02642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_137_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10232__A2 _00758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08092__I _01769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11350_ _05222_ _05441_ _05442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_137_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10301_ as2650.holding_reg\[2\] _04423_ _04436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_10_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_180_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11281_ as2650.stack\[9\]\[5\] _01934_ _01914_ as2650.stack\[8\]\[5\] as2650.stack\[10\]\[5\]
+ _01912_ _05375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_4_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10232_ _03877_ _00758_ _00926_ _02760_ _04381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XANTENNA__09925__A2 _04081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_105_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10163_ _00808_ _00608_ _04314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07436__I _01746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09689__A1 _03797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10094_ net41 _04246_ _04247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_114_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10299__A2 _02850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_142_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10797__I _04331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06911__A2 _01221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11248__A1 _05160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11727__CLK clknet_leaf_88_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10996_ _04532_ _05080_ _05095_ _03757_ _04744_ _05096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_167_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_147_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09861__A1 _04007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_163_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11617_ _05638_ _04429_ _04430_ _00756_ _05658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__11877__CLK clknet_leaf_99_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08416__A2 _02690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10223__A2 _00700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11420__A1 _02110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11548_ _05589_ _05556_ _05594_ _04298_ _05595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_183_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08931__S _03127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_171_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11479_ _02604_ _05537_ _05538_ _05539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__06442__A4 _00887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11577__B _05611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_139_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07346__I _01781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06250__I _00549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05971_ _00429_ _00430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_25_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07710_ _02122_ _02092_ _02123_ _02130_ _00037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_08690_ _00951_ _02959_ _02961_ _02817_ _02962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__07155__A2 _01454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09561__I _03724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08352__A1 _02505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07641_ _02066_ _02067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_65_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06902__A2 _01333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11239__A1 as2650.stack\[5\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11239__B2 as2650.stack\[7\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07572_ _01993_ _02000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_50_wb_clk_i clknet_4_13_0_wb_clk_i clknet_leaf_50_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08104__A1 _02394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09311_ _02631_ _03518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_59_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06523_ _00963_ _00966_ _00967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09852__A1 _03975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09852__B2 _04009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09242_ _03449_ _03450_ _03447_ _03460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_61_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06454_ _00468_ _00571_ _00897_ _00899_ _05678_ _00900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__09510__B _03640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08905__I _01309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09173_ _05765_ _03393_ _03394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09604__A1 _02844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06385_ _05696_ _00830_ _00831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_175_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08126__B _02435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08124_ _02412_ _02454_ _02460_ _02462_ _00119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06425__I _00666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11411__A1 _03555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08055_ as2650.stack\[12\]\[5\] _02396_ _02410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_174_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_134_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput17 net17 io_oeb[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__12032__CLK clknet_leaf_56_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07006_ _01133_ _01445_ _01446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput28 net28 io_out[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__09907__A2 _03788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput39 net39 io_out[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_192_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08040__B1 _02395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07256__I _01692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08591__A1 _02809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08957_ _01597_ _03119_ _03198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_4616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08796__B _03021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07908_ _02174_ _02285_ _02286_ _02295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_4649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08888_ _03077_ _03133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09471__I _00616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07146__A2 _01583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08343__A1 _02249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_99_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07839_ as2650.stack\[13\]\[9\] _02242_ _02243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__10150__A1 net92 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_99_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10850_ _00794_ _04192_ _04955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_44_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_38_wb_clk_i_I clknet_4_6_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09509_ _00572_ _02553_ _03674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10781_ _04875_ _00628_ _04888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09843__A1 _03958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08646__A2 _02913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_164_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_142_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10285__C _00911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11402_ _03542_ _05473_ _05474_ _05477_ _00382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_172_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11402__A1 _03542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06335__I _00784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09071__A2 _03257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_193_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07082__A1 _05775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11333_ _01029_ _02867_ _03679_ _00810_ _05425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_181_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11264_ _05355_ _05356_ _05357_ _05358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_140_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_140_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07909__A1 _02091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10215_ net91 _04362_ _04364_ _04365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__07909__B2 _02295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_190_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11195_ _03149_ _02833_ _05288_ _05290_ _05291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_171_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07385__A2 _01816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10146_ _03779_ _04298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_121_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_77_wb_clk_i_I clknet_4_11_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11469__A1 _00884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10077_ _04150_ _04169_ _04230_ _04231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08334__A1 _02519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08885__A2 _03108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10692__A2 _03957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_3 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_44_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_50_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10979_ net71 _05078_ _05079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_43_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06648__A1 _01080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10476__B _04588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05871__A2 _05683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06170_ _00628_ _00629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09062__A2 _03257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_1826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07073__A1 _05764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09556__I _03719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_193_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09860_ _02107_ _03959_ _04018_ _04019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08811_ _00923_ _00927_ _00931_ _03053_ _03058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XTAP_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09791_ net34 _03951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10380__A1 _01431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08742_ _02997_ _03004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05954_ _05756_ _05808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_85_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07128__A2 _00829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09291__I _03495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07804__I _02213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08673_ _02848_ _01234_ _02836_ _02940_ _02945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_26_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05885_ _05707_ _05739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10132__A1 net68 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07624_ _02050_ _02051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_26_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07555_ _01030_ _01983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09825__A1 _02613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08628__A2 _02899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_179_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06639__A1 _01061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06506_ _00949_ _00950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10435__A2 _04536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07486_ as2650.stack\[2\]\[12\] _01865_ _01872_ _01918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_39_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08635__I _02906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09225_ _03439_ _03443_ _03444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_158_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06437_ _00849_ _00883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__11061__I _05159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09428__I1 _03279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09156_ _03344_ _03373_ _03376_ _03377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__05862__A2 _05715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06368_ _00739_ _00625_ _00813_ _00814_ _00006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_175_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08107_ _02449_ _02442_ _02446_ _02450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09087_ _05758_ _01379_ _03310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_163_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06299_ _00750_ _00751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_107_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08800__A2 _02475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05994__I _05691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_190_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10833__C _00760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06811__A1 _01015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08370__I _02033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08038_ _02256_ _02397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_159_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_111_wb_clk_i_I clknet_4_3_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10000_ as2650.addr_buff\[0\] _04156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_5114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_172_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10371__A1 _03138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09989_ _02889_ _04145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_5147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07714__I net70 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output49_I net49 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11951_ _00320_ clknet_leaf_49_wb_clk_i as2650.idx_ctrl\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_4479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_177_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_84_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10902_ _04454_ _05002_ _05005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11882_ _00251_ clknet_leaf_103_wb_clk_i as2650.stack\[4\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08973__C _03127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10833_ _03639_ _01800_ _04938_ _00760_ _04939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__08619__A2 _02804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_13_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11623__A1 _02616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08545__I _00613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10764_ _04790_ _04845_ _04871_ _00732_ _04872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_164_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09292__A2 _03504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10695_ _04802_ _04803_ _04804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_40_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09419__I1 _01102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07055__A1 _01092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_153_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11316_ _05170_ _05408_ _05409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11915__CLK clknet_leaf_73_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08280__I _00873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_10_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11247_ as2650.stack\[8\]\[4\] _01961_ _05310_ as2650.stack\[11\]\[4\] _05342_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_190_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08555__A1 net94 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11178_ _05271_ _05274_ _05275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10129_ _02216_ _01609_ _04281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11574__C _03661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07624__I _02050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10114__A1 _04248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10665__A2 _01809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09979__C _03777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07530__A2 _01959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09807__A1 _00816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09807__B2 _03917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07340_ _01775_ _01776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_91_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_91_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_149_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09283__A2 _02673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07271_ _01225_ _01707_ _01708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07294__A1 net86 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11090__A2 _05188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09010_ _02302_ _02495_ _03216_ _03242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06222_ _00679_ _00680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__05844__A2 _05690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07046__A1 _01478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_1623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06153_ _00611_ _00588_ _00612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_145_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09286__I _02670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_145_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06084_ _00469_ _00542_ _00543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09912_ _03724_ _04069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10225__I _00702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07349__A2 _01740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09843_ _03958_ _02858_ _04001_ _04002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_112_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10353__A1 _03991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_154_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06986_ _01301_ _01426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09774_ _03907_ _03910_ _03934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_100_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05937_ _05789_ _05790_ _05791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_39_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08725_ _02409_ _02985_ _02988_ _02990_ _00192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_73_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_167_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11302__B1 _05157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08656_ _02135_ _02849_ _01436_ _02927_ _02928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_2329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05868_ _05720_ _05721_ _05722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_26_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07607_ _02030_ _02031_ _02034_ _02035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_54_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08587_ _02859_ _02860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_41_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11931__D _00300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05989__I _00447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10408__A2 _02573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11605__A1 _00824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07538_ as2650.stack\[9\]\[14\] _01859_ _01941_ as2650.stack\[8\]\[14\] as2650.stack\[10\]\[14\]
+ _01870_ _01968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XANTENNA__09274__A2 _03483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06088__A2 _00546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08482__B1 _01986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07469_ _01784_ _01899_ _01901_ _01902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_50_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09208_ _03385_ _03402_ _03427_ _03428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05835__A2 _05688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11938__CLK clknet_leaf_38_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10480_ _00780_ _04581_ _04593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_154_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09139_ _03357_ _03360_ _03361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_108_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07588__A2 as2650.last_intr vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_194_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10592__A1 _03914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11101_ _02811_ _00760_ _05197_ _05198_ _05199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_151_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06260__A2 _00692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11032_ _05130_ _05131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_2_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10344__A1 _00811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10344__B2 _00825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06012__A2 _00470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06563__A3 _01003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07760__A2 _02172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08984__B _02501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11934_ _00303_ clknet_leaf_61_wb_clk_i net39 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10647__A2 _04755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_146_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07512__A2 _01940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11865_ _00234_ clknet_leaf_29_wb_clk_i as2650.r123_2\[0\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_17_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_177_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_107_wb_clk_i clknet_4_3_0_wb_clk_i clknet_leaf_107_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_60_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10816_ _02194_ _04914_ _04922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_18_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11796_ _00179_ clknet_leaf_124_wb_clk_i as2650.stack\[15\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_158_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09265__A2 _03443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07276__A1 _00605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10747_ _04023_ _04801_ _04855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_70_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10678_ _04532_ _04748_ _04773_ _04787_ _04744_ _04788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_185_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07028__A1 _01466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_182_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07579__A2 _00626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07619__I _02046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08776__A1 _02976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10583__A1 _01776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08240__A3 _02548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06251__A2 _00545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08528__A1 as2650.stack\[13\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08528__B2 as2650.stack\[12\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11585__B _05629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06840_ _01016_ _00977_ _01282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__06003__A2 _00461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10886__A2 _04979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07354__I _01789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06771_ _05814_ _01134_ _01110_ _01212_ _01213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_42_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08510_ as2650.stack\[7\]\[6\] _02782_ _01780_ as2650.stack\[6\]\[6\] _02783_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_48_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09490_ _00504_ _03657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_110_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08441_ _02706_ _02717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_1_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08372_ _02665_ _02666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_189_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09256__A2 _03342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07323_ as2650.stack\[5\]\[8\] _01753_ _01758_ as2650.stack\[4\]\[8\] _01759_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_32_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_177_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07254_ _01257_ _01690_ _01691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_140_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09008__A2 _03233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_191_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06205_ as2650.ins_reg\[2\] _00447_ _00664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_10_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07185_ _01225_ _01622_ _01623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07529__I _01874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06136_ _00589_ _05787_ _00595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__06433__I _00878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10574__A1 as2650.stack\[2\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10574__B2 as2650.stack\[0\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06067_ _00512_ _00522_ _00525_ _00526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__08519__A1 _02789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07990__A2 _02222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10326__A1 _04454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09192__A1 _03395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11926__D _00295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09826_ _03978_ _01444_ _03985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_100_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09757_ _03909_ _03918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_58_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06969_ _01398_ _01406_ _01408_ _01409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
Xclkbuf_leaf_5_wb_clk_i clknet_4_1_0_wb_clk_i clknet_leaf_5_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_55_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08708_ _02971_ _02978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09688_ _03849_ _03850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_15_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08639_ as2650.stack\[5\]\[7\] _01790_ _01794_ as2650.stack\[4\]\[7\] _02911_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_128_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11650_ _00033_ clknet_leaf_134_wb_clk_i as2650.stack\[13\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_184_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06608__I _01051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_19_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11760__CLK clknet_leaf_81_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_3_0_0_wb_clk_i_I clknet_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07258__A1 _01601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10601_ _04454_ _04702_ _04712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07258__B2 _01319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11581_ _02956_ _02609_ _05626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xfanout85 net29 net85 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_195_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10532_ _04404_ _04645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_168_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08823__I _03066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10801__A2 _04878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_167_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_109_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06481__A2 _00484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10463_ _04554_ _04575_ _04576_ _04577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_136_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08758__A1 _02409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09955__B1 _04111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06343__I _00792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10394_ _02837_ _04484_ _04510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10565__A1 _04226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06233__A2 _00690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07430__A1 as2650.stack\[3\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_150_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10317__A1 _05674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11015_ _00864_ _05113_ _02806_ _05114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_104_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08930__A1 _01429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_92_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09486__A2 _00504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08289__A3 _02597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11917_ _00286_ clknet_leaf_73_wb_clk_i as2650.stack\[5\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11848_ _00008_ clknet_leaf_48_wb_clk_i as2650.cycle\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_53_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09238__A2 _03338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11779_ _00162_ clknet_leaf_93_wb_clk_i as2650.stack\[3\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_144_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08997__A1 _03037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10484__B net56 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_75_wb_clk_i clknet_4_11_0_wb_clk_i clknet_leaf_75_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_103_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11348__A3 _05439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09410__A2 _02514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06224__A2 _00681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08990_ _02368_ _02500_ _03227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09564__I _03727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_114_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07941_ _02280_ _02317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10308__A1 as2650.holding_reg\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05983__A1 _05704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11633__CLK clknet_leaf_27_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_190_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10859__A2 _04961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07872_ _02227_ _02263_ _02264_ _02265_ _00064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_131_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08921__A1 _03110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09611_ _03759_ _03770_ _03772_ _03773_ _03774_ _03775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_06823_ _05766_ _01265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_28_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06754_ _01115_ _01197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_110_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09542_ _00735_ _00729_ _03704_ _03705_ _03706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_37_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09477__A2 _00772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11783__CLK clknet_leaf_85_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06685_ _00637_ _00979_ _01128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09473_ _00622_ _00687_ _03640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07488__B2 as2650.stack\[8\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11284__A2 _05377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08424_ _02686_ _02700_ _02701_ _02704_ _00177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_93_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06160__A1 _00586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06428__I _00873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08355_ _02513_ _02646_ _02652_ _02654_ _00158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_75_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06872__B _01027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08988__A1 _02364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07306_ net48 _01742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_149_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08286_ _00597_ _00603_ _02573_ _02595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_20_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10795__A1 _03824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08452__A3 _02724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07237_ _01669_ _01674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_165_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06463__A2 _00586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07660__A1 _01905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_121_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07259__I _01695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_118_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07168_ _05801_ _01605_ _01606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_195_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10547__A1 _04200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09401__A2 _03575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06215__A2 _00661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06119_ _00480_ _00457_ _00578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_132_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07099_ _01393_ _01201_ _01523_ _01537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__07412__B2 _01846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09474__I _02823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_182_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08311__C _02619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08912__A1 _01306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09809_ _03958_ _03959_ _03967_ _03968_ _03969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_19_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06774__I0 as2650.r123\[0\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06923__B1 _01363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08818__I _03064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output31_I net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07722__I _01782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09468__A2 _03627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_56_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08140__A2 _02475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11702_ _00085_ clknet_leaf_116_wb_clk_i as2650.stack\[10\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06151__A1 _00606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11633_ _00016_ clknet_leaf_27_wb_clk_i as2650.r123\[1\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08979__A1 _02648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08553__I _01610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_180_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_54_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11564_ _02076_ _05597_ _05606_ _05609_ _05610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_156_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10786__A1 _04883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06454__A2 _00571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10515_ as2650.stack\[3\]\[1\] _01835_ _02909_ as2650.stack\[2\]\[1\] _04628_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_11495_ _05549_ _00403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07169__I net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10446_ _02037_ _00513_ _04560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_100_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_170_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07403__A1 as2650.stack\[10\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10377_ _03267_ _04490_ _04496_ _04497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_151_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09384__I _03574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07954__A2 _02319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05965__A1 _05789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12047_ _00416_ clknet_4_4_0_wb_clk_i net50 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_117_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08903__A1 _01156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08903__B2 _01318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_122_wb_clk_i clknet_4_0_0_wb_clk_i clknet_leaf_122_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_92_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06390__A1 _00511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09459__A2 _03627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08667__B1 _01042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11266__A2 _02960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08667__C2 _02854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_178_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06470_ _00508_ _00599_ _00912_ _00915_ _00891_ _00916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_33_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11018__A2 _04319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09559__I _03722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08140_ as2650.stack\[8\]\[9\] _02475_ _02476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_33_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06445__A2 _00545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08071_ _02422_ _02423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07642__A1 as2650.stack\[13\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_174_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07079__I _01517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07022_ _05744_ _05748_ _01461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09395__A1 _02167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07807__I net67 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07945__A2 _02319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06711__I _01132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08973_ _01693_ _03071_ _03212_ _03127_ _03213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_103_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07924_ _02304_ _02197_ _02305_ _02306_ _00075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_4809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_57_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07855_ as2650.stack\[12\]\[8\] _02251_ _02253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__10701__A1 _02952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06806_ _01082_ _01238_ _01244_ _01077_ _01247_ _01248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
XFILLER_99_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07786_ _02029_ _02198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_84_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09525_ _00772_ _00784_ _01712_ _02580_ _03689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_06737_ _01179_ _01180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11257__A2 _01501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11064__I _01941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xclkbuf_3_5_0_wb_clk_i clknet_0_wb_clk_i clknet_3_5_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_73_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_06668_ _01111_ _01112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_40_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09456_ _02534_ _03627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_94_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09870__A2 _01457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__11009__A2 _00599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08407_ _02693_ _02694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_51_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06599_ _01042_ _01043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_123_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09387_ as2650.stack\[6\]\[0\] _03577_ _03578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_178_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09469__I net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_184_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08338_ _02521_ _02639_ _02640_ _02641_ _00154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__08425__A3 _02664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11679__CLK clknet_leaf_131_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08269_ _00734_ _01037_ _02562_ _02577_ _02578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_126_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10232__A3 _00926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10300_ _04433_ _04434_ _04435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_137_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11280_ as2650.stack\[11\]\[5\] _02002_ _05374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_152_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_180_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10231_ _00564_ _00556_ _04379_ _03644_ _04380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_49_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07717__I _02136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07936__A2 _02160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output79_I net79 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06621__I _05734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10162_ _00782_ _02737_ _03678_ _04313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_120_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09138__A1 _05764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_67_wb_clk_i_I clknet_4_12_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10093_ _04209_ _04210_ _04246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_120_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08649__B1 _01814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10995_ _01974_ _04995_ _05093_ _05094_ _05095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_188_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09310__A1 _03050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_95_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09861__A2 _03724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07872__A1 _02227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09379__I _02121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11616_ _04460_ _05575_ _05647_ _05657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_30_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10759__A1 _02351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06427__A2 _00872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__11420__A2 _05462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11547_ _02027_ _05579_ _05593_ _05594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_156_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06978__A3 _01417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11478_ _02565_ _04523_ _05538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__09377__A1 _03239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10429_ as2650.stack\[3\]\[0\] _04536_ _04542_ as2650.stack\[2\]\[0\] _04543_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_140_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11184__A1 _03974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07627__I net56 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10481__C _02334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07927__A2 _02207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10931__A1 _05031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09129__A1 _03327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05970_ _05779_ _00429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_140_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_66_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07640_ _02065_ _02066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07571_ _01991_ _01999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_53_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11239__A2 _05302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08104__A2 _02436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09301__A1 _03040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06522_ _00965_ _00966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09310_ _03050_ _03508_ _03516_ _03517_ _00250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_165_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07312__B1 _01747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_181_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09852__A2 _03742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10998__A1 _00799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09241_ _03434_ _03457_ _03458_ _03459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_146_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06453_ _00500_ _00898_ _00899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_107_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07863__A1 _02207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_194_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09289__I _02665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_90_wb_clk_i clknet_4_8_0_wb_clk_i clknet_leaf_90_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_09172_ _01649_ _03393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06384_ _00829_ _00830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_119_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08123_ _02461_ _02425_ _02435_ _02462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__07615__A1 _01100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07030__C _01468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11411__A2 _05473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08054_ _02101_ _02409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_179_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11971__CLK clknet_leaf_39_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07005_ _01444_ _01445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09368__A1 as2650.stack\[3\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_101_wb_clk_i_I clknet_4_3_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput18 net18 io_oeb[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput29 net29 io_out[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_162_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11175__A1 as2650.stack\[9\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08040__A1 _02394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10922__A1 _04999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_89_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08956_ _02835_ _03133_ _03196_ _03075_ _03197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_4606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07907_ as2650.stack\[10\]\[4\] _02293_ _02294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_4639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11478__A2 _04523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08887_ _01262_ _03075_ _03132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_3905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_56_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09540__A1 _03702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08343__A2 _02630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07838_ _02035_ _02242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_57_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06354__A1 _00713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_183_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07769_ _02113_ _02172_ _02180_ _02182_ _00044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_25_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09508_ _02581_ _03673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_169_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06106__A1 _00536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10780_ _03921_ _00895_ _04608_ _04886_ _04887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_53_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09843__A2 _02858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10989__A1 _04897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09439_ _02003_ _03024_ _03218_ _03614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XPHY_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_157_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10566__C _00521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_185_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11401_ as2650.stack\[9\]\[0\] _05476_ _05468_ _05477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_122_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06409__A2 _00767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11402__A2 _05473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08831__I _03077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11332_ _05142_ _00759_ _05423_ _05424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_180_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09359__A1 as2650.stack\[3\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11263_ _05249_ _01518_ _05357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_137_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07909__A2 _02292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10214_ _04363_ _04364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08031__A1 as2650.stack\[12\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06351__I _00799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11194_ _03148_ _02815_ _05249_ _05289_ _05241_ _05290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_133_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10913__A1 _04604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10145_ _02225_ _04111_ _04296_ _00452_ _04297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__07891__B _02281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11469__A2 _04349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10076_ net87 _02193_ _04229_ _04230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_48_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09531__A1 _00832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_4_10_0_wb_clk_i_I clknet_3_5_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10677__B1 _04786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09531__B2 _00778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10692__A3 _02080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_189_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10429__B1 _04542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08098__A1 _02276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10978_ _05055_ _05031_ _05078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_147_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_71_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06648__A2 _01091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07845__A1 as2650.stack\[13\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06526__I _00946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11994__CLK clknet_4_5_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_30_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_141_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08270__A1 _02571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_1849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11157__A1 _02841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08022__A1 as2650.stack\[14\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08897__B _03141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08810_ _03056_ _03057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09770__A1 _03886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09790_ _03941_ _03942_ _03949_ _03950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_119_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08741_ _02976_ _02700_ _03003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05953_ _05805_ _05806_ _05807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05884_ as2650.r123\[1\]\[5\] as2650.r123\[0\]\[5\] as2650.r123_2\[1\]\[5\] as2650.r123_2\[0\]\[5\]
+ _05684_ _05736_ _05738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_08672_ _01141_ _01034_ _01297_ _02853_ _02944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_27_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08188__I _02510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10132__A2 _02940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07533__B1 _01962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07623_ _02049_ _02050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_53_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08089__A1 _02329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07554_ _01979_ _01910_ _01982_ _00029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_74_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09825__A2 _03887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06505_ _00948_ _00449_ _00949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_34_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07485_ as2650.stack\[3\]\[12\] _01862_ _01863_ as2650.stack\[0\]\[12\] _01753_ as2650.stack\[1\]\[12\]
+ _01917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_22_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09224_ _03441_ _03442_ _03443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_166_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06436_ _00881_ _00882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06436__I _00881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_3_5_0_wb_clk_i_I clknet_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09589__A1 _03749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09155_ _03346_ _03372_ _03376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06367_ _00720_ _00691_ _00814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_124_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08106_ _02073_ _02449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_87_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_174_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09086_ _01635_ _01644_ _03309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_162_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06298_ _00747_ _05678_ _00749_ _00750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_174_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11929__D _00298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08037_ _02389_ _02396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06811__A2 _00432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11717__CLK clknet_leaf_134_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06171__I _00629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10746__I1 _04853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_137_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09761__A1 _03886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_5115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09988_ _00633_ _04143_ _04144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_5137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08939_ _02933_ _03114_ _03115_ _03180_ _03181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_131_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11517__I _02746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09513__A1 _02823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10421__I _04534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11950_ _00319_ clknet_leaf_49_wb_clk_i as2650.idx_ctrl\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_4469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06327__A1 _00564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10901_ _03820_ _04262_ _05003_ _05004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_57_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11881_ _00250_ clknet_leaf_97_wb_clk_i as2650.stack\[2\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_45_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10832_ _03639_ _04934_ _04938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08826__I _03072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10763_ _04869_ _04870_ _04871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_158_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10694_ _02094_ _04704_ _02107_ _04803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_142_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11387__A1 _02678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_154_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09657__I _02952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08561__I _01602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08252__A1 _00605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_181_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11839__D _00222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_177_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11315_ _05404_ _05407_ _05408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_126_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11139__A1 _03974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05861__I0 as2650.r123\[1\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06081__I _00531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08004__A1 as2650.stack\[14\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11246_ as2650.stack\[10\]\[4\] _05225_ _05178_ as2650.stack\[9\]\[4\] _05341_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_122_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09752__A1 _00731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08555__A2 _02826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06566__A1 _01008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11177_ _05160_ _05272_ _05273_ _05274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_110_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09392__I _02511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07905__I _02280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10128_ _04216_ _04249_ _04280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_5660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09504__A1 net24 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_5693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10059_ _02204_ _01611_ _04213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_4970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_29_wb_clk_i clknet_4_7_0_wb_clk_i clknet_leaf_29_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_36_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_169_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_90_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12022__CLK clknet_leaf_38_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09268__B1 _03340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09807__A2 _03961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07640__I _02065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07818__A1 _02223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07818__B2 _02225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07270_ _01226_ _01686_ _01706_ _01707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_149_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06256__I _00711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07294__A2 _01729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05924__S0 as2650.ins_reg\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06221_ _00523_ _00679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_31_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06152_ _00595_ _00611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_89_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07046__A2 _00667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10050__A1 _04200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06083_ as2650.prefixed _05699_ _00542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_160_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_1679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09911_ _04067_ _04068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_67_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09043__I0 _03270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09743__A1 _03811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09842_ _03933_ _03935_ _04001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_112_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07815__I _01380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08420__B _02701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11550__A1 _02027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09773_ _03932_ _03933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_112_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06985_ _01308_ _05810_ _01425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_101_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08724_ _02989_ _02712_ _02969_ _02990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_160_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05936_ _05779_ _05790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_113_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11302__A1 as2650.stack\[6\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11302__B2 as2650.stack\[4\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08655_ net74 _02927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_26_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05867_ as2650.r123\[2\]\[7\] as2650.r123_2\[2\]\[7\] _05713_ _05721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_82_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07606_ _02033_ _02034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_1618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08586_ _02858_ _02859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_82_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07550__I as2650.r123\[0\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_165_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07537_ _01965_ _01966_ _01799_ _01967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__11605__A2 _02903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_180_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11072__I _01812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06166__I _00547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_167_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07468_ as2650.stack\[13\]\[11\] _01900_ _01879_ as2650.stack\[12\]\[11\] _01901_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08482__B2 _00606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_194_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09207_ _03387_ _03401_ _03427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06419_ _00864_ _00865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_195_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07399_ _01831_ _01833_ _01777_ _01834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09138_ _05764_ _01542_ _03360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07037__A2 _01471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08234__A1 _02525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10416__I _04529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07588__A3 net75 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09069_ _03284_ _03292_ _03293_ _00233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_151_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10592__A2 _04646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_162_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11100_ _03148_ _02833_ _05198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_150_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10860__B _04374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11031_ _00851_ _00872_ _00845_ _05130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_172_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10344__A2 _00751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output61_I net61 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11541__A1 _04460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_134_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06563__A4 _01006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11933_ _00302_ clknet_leaf_61_wb_clk_i net38 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_185_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11864_ _00233_ clknet_leaf_29_wb_clk_i as2650.r123_2\[0\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10815_ _00809_ _04152_ _04920_ _04921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_57_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11795_ _00178_ clknet_leaf_123_wb_clk_i as2650.stack\[15\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09265__A3 _03470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06076__I net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10746_ _04846_ _04853_ _04608_ _04854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07276__A2 _01711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10280__A1 _04415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10677_ _04535_ _04749_ _04786_ _04742_ _04640_ _04787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_126_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08225__A1 as2650.stack\[5\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10032__A1 _04186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10032__B2 _04181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08776__A2 _03029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06787__A1 as2650.holding_reg\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08528__A2 _02785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11229_ _02724_ _04786_ _05323_ _05134_ _05324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_136_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06539__A1 _00709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11585__C _00756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11532__A1 _01986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07635__I _02024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06770_ _01199_ _01212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_97_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_95_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09850__I _00698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_110_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08440_ _02678_ _02707_ _02711_ _02716_ _00181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__08700__A2 _02001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08371_ _02186_ _02649_ _02664_ _02665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_149_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11599__A1 _03972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07322_ _01757_ _01758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07267__A2 _01696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10271__A1 _04409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06475__B1 _00890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07253_ _01600_ _01689_ _01690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_143_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09297__I _02670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_192_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06204_ _00589_ _00663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07184_ _01226_ _01589_ _01621_ _01622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_121_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08216__A1 as2650.stack\[5\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10023__A1 _04156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09964__A1 _00961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06135_ _00588_ _00593_ _00594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__10236__I _04384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_191_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06778__A1 _01020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10574__A2 _04681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06066_ _00523_ _00524_ _00525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09716__A1 _03665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_120_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07545__I _01598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10326__A2 _00783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08150__B _02481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11523__A1 _04437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09192__A2 _03399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09825_ _02613_ _03887_ _01005_ _03984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_115_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09756_ _03817_ _03917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_58_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06968_ _01180_ _01188_ _01407_ _01408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09760__I _01697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_27_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08707_ _02976_ _02717_ _02977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05919_ as2650.ins_reg\[4\] _05772_ _05773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09687_ _00980_ _03849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06899_ _01335_ _01338_ _01339_ _01340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_54_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08638_ as2650.stack\[7\]\[7\] _02908_ _02909_ as2650.stack\[6\]\[7\] _02910_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_54_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11905__CLK clknet_leaf_72_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11016__B _05114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08569_ _02841_ _02842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_180_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10600_ _03914_ _03734_ _04710_ _04711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_106_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07258__A2 _01017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08455__A1 _02723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11580_ _01327_ _01416_ _01421_ _05625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_23_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_126_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout86 net59 net86 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10262__A1 as2650.last_intr vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10531_ _04533_ _04582_ _04619_ _04641_ _04643_ _04644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_52_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10462_ _03749_ _04556_ _03738_ _00672_ _04576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_108_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09955__A1 _03830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08758__A2 _03011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11211__B1 _05172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10146__I _03779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09955__B2 _02126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10393_ _04489_ _04508_ _04509_ _00341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__06769__A1 _01210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10565__A2 _04676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07430__A2 _01862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09707__A1 _00630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07455__I as2650.r123\[0\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10317__A2 _04399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11514__A1 _05561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11014_ _03650_ _01131_ _05110_ _05112_ _00555_ _05113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_81_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_49_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06941__A1 _05776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_77_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_189_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11278__B1 _01936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10749__C _02901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11916_ _00285_ clknet_leaf_94_wb_clk_i as2650.stack\[5\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07497__A2 _01926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08694__A1 _02843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11847_ _00007_ clknet_leaf_47_wb_clk_i as2650.cycle\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_127_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08446__A1 _02684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11778_ _00161_ clknet_leaf_93_wb_clk_i as2650.stack\[3\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_13_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11450__B1 _05513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10729_ _04535_ _04793_ _04837_ _04742_ _04062_ _04838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_105_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06534__I _00977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08749__A2 _02998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09845__I _03776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_4_7_0_wb_clk_i clknet_3_3_0_wb_clk_i clknet_4_7_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_142_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_102_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07940_ as2650.stack\[10\]\[8\] _02297_ _02316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_69_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10308__A2 _04423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11505__A1 _04437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05983__A2 _05693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_155_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07871_ as2650.stack\[12\]\[12\] _02260_ _02265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_116_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10859__A3 _04962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09610_ _00551_ _03774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08921__A2 _03162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06822_ _01051_ _01264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_55_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09580__I _03743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09541_ _00891_ _02005_ _02572_ _03705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_06753_ _01164_ _01195_ _01000_ _01196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_clkbuf_leaf_18_wb_clk_i_I clknet_4_5_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07488__A2 _01869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08196__I _02506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09472_ _03638_ _03639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_168_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06684_ _01125_ _01126_ _01127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08685__A1 _02951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10492__A1 _04604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08423_ as2650.stack\[1\]\[14\] _02689_ _02704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_63_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_145_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08354_ as2650.stack\[3\]\[9\] _02653_ _02654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_149_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10675__B _04784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10244__A1 _01274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07305_ net86 _01741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__08988__A2 _03222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08285_ _02592_ _02593_ _02567_ _01038_ _02594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_20_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06999__A1 _01433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10795__A2 _04901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07236_ _01671_ _01672_ _01673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_30_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07167_ _00942_ _01604_ _01605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_173_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10547__A2 _03960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09755__I _03915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06118_ _00523_ _00574_ _00576_ _00577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_136_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06215__A3 _00671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07098_ _01509_ _01534_ _01535_ _01536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_161_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06049_ _00506_ _00507_ _00508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_57_wb_clk_i_I clknet_4_15_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05974__A2 _00431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07176__A1 _01599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09808_ _03878_ _03968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_60_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09490__I _00504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06923__B2 _01020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09739_ _03894_ _03898_ _03899_ _03900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_74_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_4_15_0_wb_clk_i_I clknet_3_7_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08676__A1 _01466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output24_I net24 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11701_ _00084_ clknet_leaf_116_wb_clk_i as2650.stack\[10\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06151__A2 _00608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11632_ _00015_ clknet_leaf_36_wb_clk_i as2650.r123\[1\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_126_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08979__A2 _02000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11563_ _00471_ _02757_ _02734_ _05608_ _05609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_168_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07100__A1 _01393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10514_ as2650.stack\[1\]\[1\] _01829_ _01826_ as2650.stack\[0\]\[1\] _04627_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_128_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11494_ as2650.r123\[3\]\[4\] _05549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_96_wb_clk_i_I clknet_4_9_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10445_ _04418_ _04558_ _04559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_152_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07403__A2 _01812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10376_ _03148_ _04491_ _04496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11847__D _00007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12046_ _00415_ clknet_leaf_16_wb_clk_i net51 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_49_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_172_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08903__A2 _01298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06390__A2 _00835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07134__B _01571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_opt_2_0_wb_clk_i clknet_4_10_0_wb_clk_i clknet_opt_2_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_52_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08667__A1 _05687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08667__B2 _01030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_178_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10226__A1 _00880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08070_ _02153_ _01989_ _01995_ _02422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__07642__A2 _02025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07021_ _01390_ _01460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_134_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09575__I _01042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10942__C _05043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08972_ _03073_ _03210_ _03211_ _03093_ _03212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_114_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_9_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07923_ _02157_ _02306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11750__CLK clknet_leaf_113_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_190_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10450__S _04563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07854_ _02251_ _02252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08919__I _03103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06905__A1 _00884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06805_ _01086_ _01246_ _01236_ _01088_ _01165_ _01247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_84_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07785_ _02196_ _02197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_71_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10389__C _04506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09524_ _00616_ _02593_ _03688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06736_ _01178_ _01173_ _01174_ _01179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__06439__I _00884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10465__A1 _03916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09455_ _03558_ _03613_ _03625_ _03626_ _00286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06667_ _01110_ _01111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_25_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_51_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08406_ _02692_ _02693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_169_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_130_wb_clk_i_I clknet_4_0_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09386_ _03576_ _03577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_75_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06598_ _01041_ _01042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_40_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10217__A1 net91 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08337_ as2650.stack\[4\]\[12\] _02636_ _02641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09083__A1 _01547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06174__I _00632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11013__C _01130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08830__A1 _01026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08268_ _02012_ _00841_ _02577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_137_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10232__A4 _02760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07219_ _01631_ _01655_ _01656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_152_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08199_ _02219_ _02519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10230_ _02806_ _02747_ _04379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_134_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10161_ _00546_ _04311_ _04312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_175_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10940__A2 _05041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09138__A2 _01542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10092_ _04129_ _04243_ _04244_ _04024_ _04245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__07149__A1 _01341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08897__A1 _03122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_47_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06349__I _00448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09846__B1 _04003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08649__B2 as2650.stack\[13\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10994_ _04535_ _05080_ _05094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_15_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09310__A2 _03508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06793__B _01232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08564__I _02836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07872__A2 _02263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11615_ _02077_ _05653_ _05656_ _00712_ _00416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__09074__A1 _00514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_15_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10759__A2 _04845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11546_ _05590_ _05565_ _05592_ _02621_ _05566_ _05593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__08821__A1 _00921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11477_ _04346_ _05527_ _05528_ _05536_ _05537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_137_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10762__C _04062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09377__A2 _02653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10428_ _01743_ _04542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_139_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11184__A2 _05280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10359_ _04480_ _04481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_139_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_191_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06968__B _01407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12029_ _00398_ clknet_4_4_0_wb_clk_i net48 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_65_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07643__I net89 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10695__A1 _04802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07570_ _01997_ _01998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_47_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10002__C _03925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06521_ _00964_ _00926_ _00965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09301__A2 _03508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07312__A1 as2650.stack\[7\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07312__B2 as2650.stack\[6\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10998__A2 _05671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09240_ _03435_ _03452_ _03458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__10937__C _04891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06452_ _00589_ _00587_ _00898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08474__I _00703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07863__A2 _02252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06910__I1 _01350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09171_ _03388_ _03391_ _03392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_33_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09065__A1 _01975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06383_ _00828_ _00829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__10509__I _04621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_147_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_119_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08122_ _02118_ _02461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_174_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08053_ _02405_ _02406_ _02407_ _02408_ _00102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_116_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_176_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07004_ _01316_ _01424_ _01425_ _01318_ _01443_ _01444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_116_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput19 net19 io_oeb[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_190_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11175__A2 _05266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08955_ _03112_ _03195_ _03196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08591__A3 _02843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_102_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07906_ _02273_ _02293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_57_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08886_ _03110_ _03129_ _03131_ _00212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_4629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10686__A1 _01464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_56_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07837_ _02239_ _02197_ _02240_ _02241_ _00053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_3939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11075__I _05164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06169__I _00627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07768_ _02181_ _02178_ _02140_ _02182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_56_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09507_ _00483_ _02554_ _03672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__10438__A1 _01775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06719_ _01154_ _01161_ _01162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_25_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06106__A2 _00564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07699_ _02113_ _02092_ _02114_ _02120_ _00036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XPHY_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10989__A2 _05080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10847__C _04326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_188_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08384__I _02665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09438_ _03612_ _03613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_125_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_157_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_184_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08317__C _02625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09369_ _02456_ _03548_ _03553_ _03564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__10419__I _04532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11400_ _05475_ _05476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_123_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11796__CLK clknet_leaf_124_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08803__A1 _02381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_166_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11331_ _02817_ _02961_ _05417_ _05422_ _05423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_115_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06290__A1 _00739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11262_ _03149_ _02814_ _05356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_49_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11166__A2 _05262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10213_ _00702_ _04363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_121_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11193_ _01363_ _05289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__08031__A2 _02390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06042__A1 _00500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10913__A2 _05004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10144_ _00673_ _04290_ _04294_ _04295_ _04296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_95_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10075_ _04136_ _04229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_23_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11469__A3 _05062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09531__A2 _02567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07542__A1 _01766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10692__A4 _04653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10429__A1 as2650.stack\[3\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_62_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10429__B2 as2650.stack\[2\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_186_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09611__C _03774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09295__A1 _03231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10977_ _02235_ _05077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_95_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07845__A2 _02242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_189_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_148_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_175_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09047__A1 _03273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10329__I _04456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06805__B1 _01236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10601__A1 _04454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_1817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11529_ _02648_ _02152_ _05577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_195_1828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08270__A2 _02573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11157__A2 _03815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08022__A2 _02360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_84_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09770__A2 _03837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08740_ _02384_ _02996_ _02999_ _03002_ _00195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05952_ _05745_ _05761_ _05762_ _05708_ _05806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07373__I _01196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10668__A1 as2650.stack\[3\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08671_ _02939_ _02941_ _02942_ _02943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_6_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05883_ as2650.r123\[2\]\[5\] as2650.r123_2\[2\]\[5\] _05736_ _05737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_27_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07533__A1 as2650.stack\[5\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07533__B2 as2650.stack\[4\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07622_ net79 _02049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_93_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07553_ _01707_ _01911_ _01718_ _01981_ _01982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_179_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08089__A2 _02430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06504_ _00487_ _00948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11093__A1 net79 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06639__A3 _01068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07484_ _01735_ _01913_ _01915_ _01916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_179_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09223_ _05724_ _01518_ _03442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05847__A1 _05691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10239__I _04385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06435_ _00880_ _00881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09154_ _03129_ _03298_ _03375_ _00236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09589__A2 _03752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06366_ _00811_ _00717_ _00812_ _00639_ _00813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_108_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08105_ as2650.stack\[0\]\[2\] _02440_ _02448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09085_ _03306_ _03307_ _03308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06297_ _00748_ _00749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_68_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06272__A1 _00625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08036_ _02060_ _02263_ _02395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_123_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_157_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_115_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06024__A1 _00478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09761__A2 _03921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_192_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09987_ _04137_ _04141_ _04143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_118_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07772__A1 _02184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_5149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08938_ _05804_ _03082_ _03180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__10702__I _03750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08379__I _02206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_170_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10659__A1 _02858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09513__A2 _02568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08869_ _00609_ _03055_ _03115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_3714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07524__A1 _01954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06327__A2 _00690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11320__A2 _05412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10900_ _04999_ _00809_ _05003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_44_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_17_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11880_ _00249_ clknet_leaf_98_wb_clk_i as2650.stack\[2\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_189_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10831_ _00452_ _04928_ _04933_ _04936_ _04937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XANTENNA__09277__A1 _03475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10762_ _04742_ _02804_ _04845_ _04534_ _04062_ _04870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_13_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10831__A1 _00452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10693_ _00444_ _04802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_41_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11387__A2 _05457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08252__A2 _00798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11314_ _05177_ _05405_ _05406_ _05407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_180_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06362__I _00808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11139__A2 _05236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05861__I1 as2650.r123\[0\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11245_ _05338_ _05339_ _05340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09201__A1 _05743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08004__A2 _02360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05907__S _05736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09752__A2 _03782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11176_ as2650.stack\[8\]\[2\] _01914_ _01937_ as2650.stack\[11\]\[2\] as2650.stack\[10\]\[2\]
+ _01933_ _05273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_68_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06566__A2 _01009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11855__D _00002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10127_ _03759_ _04276_ _04278_ _03772_ _03774_ _04279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__10612__I _00894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09504__A2 _03669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10058_ _00718_ _04208_ _04211_ _03995_ _04004_ _04212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_57_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07921__I _02160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__11961__CLK clknet_leaf_15_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09268__A1 _03202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_69_wb_clk_i clknet_4_9_0_wb_clk_i clknet_leaf_69_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_16_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10822__A1 _04879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06220_ _00677_ _00678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_31_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09848__I net61 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08752__I _02693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_89_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06151_ _00606_ _00608_ _00585_ _00609_ _00610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_121_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06254__A1 _00694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_176_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06082_ _00540_ as2650.cycle\[11\] _00541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09910_ _03719_ _04067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06006__A1 _05700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10950__C _00882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09841_ _03999_ _04000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10889__A1 _04879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09743__A2 _03903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10889__B2 _04771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_119_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07754__A1 _02170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09772_ _02093_ net12 _03932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__08199__I _02219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06984_ _01390_ _01423_ _01424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08723_ _02109_ _02989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05935_ _05787_ _05788_ _05789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_80_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08654_ _00843_ _01090_ _00493_ _00464_ _02926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XTAP_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05866_ _05719_ _05720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_54_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10510__B1 _01790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07831__I _02236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07605_ _02019_ _02020_ _02032_ _02033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_148_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08585_ _01436_ _02858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_26_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10397__C _04506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07536_ as2650.stack\[2\]\[14\] _01944_ _01735_ _01966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__06447__I _00576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11605__A3 _02860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10813__A1 _04654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07467_ _01815_ _01900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_195_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08482__A2 _00899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09206_ _03390_ _03425_ _03426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_108_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06418_ _00863_ _00864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_183_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07398_ as2650.stack\[3\]\[9\] _01832_ _01788_ _01833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_148_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09137_ _03356_ _03324_ _03358_ _03359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_194_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06349_ _00448_ _00798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_120_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_175_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10577__B1 _01794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09068_ as2650.r123_2\[0\]\[6\] _03259_ _03293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_11_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_136_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07993__A1 as2650.stack\[14\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08019_ _02113_ _02373_ _02379_ _02380_ _00096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__11834__CLK clknet_leaf_32_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11030_ _05103_ _05129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_1_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11541__A2 _05575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output54_I net54 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11984__CLK clknet_leaf_77_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_4245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_134_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09498__A1 _03636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11932_ _00301_ clknet_leaf_61_wb_clk_i net37 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_4289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07741__I _02155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11863_ _00232_ clknet_leaf_29_wb_clk_i as2650.r123_2\[0\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10814_ _04913_ _04077_ _04920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_96_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06357__I _00804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11794_ _00177_ clknet_leaf_86_wb_clk_i as2650.stack\[1\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_158_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10804__A1 as2650.ivec\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10745_ _04025_ _04009_ _04850_ _04852_ _04853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__10804__B2 _04878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09670__A1 _03814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08572__I _02844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10676_ _04776_ _04779_ _04785_ _01844_ _04786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_173_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08225__A2 _02538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10032__A2 _00682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_177_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07984__A1 _02347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10583__A3 _04694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_116_wb_clk_i clknet_4_2_0_wb_clk_i clknet_leaf_116_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_107_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_153_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09186__B1 _03406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06820__I _01210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11228_ _00955_ _05131_ _05322_ _05323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_122_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06539__A2 _00642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11532__A2 _05177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11159_ as2650.stack\[4\]\[2\] _05210_ _05256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_190_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_191_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09489__A1 _02566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11296__A1 _01599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11296__B2 _02234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07651__I _01028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08700__A3 _02143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11048__A1 _05128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08370_ _02033_ _02664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_56_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07321_ _01756_ _01757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09578__I _03741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06475__A1 _00452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07252_ _01451_ _01308_ _01461_ _01423_ _01689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_143_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06475__B2 _05674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_164_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06203_ _00486_ _00662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__11122__B _05152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07183_ _01055_ _01617_ _01620_ _01293_ _01621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__11857__CLK clknet_4_12_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08216__A2 _02530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09413__A1 _02129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06227__A1 _00448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10023__A2 _04118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06134_ _00590_ _00592_ _00593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__11220__A1 _05264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_160_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06778__A2 _01219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07975__A1 _00811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06065_ _00487_ _00484_ _00524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_105_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_47_wb_clk_i_I clknet_4_13_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09716__A2 _03877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10326__A3 _00786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11523__A2 _05570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09824_ _03803_ _03982_ _03983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06967_ _01245_ _01236_ _01334_ _01407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09755_ _03915_ _03916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_104_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05918_ as2650.alu_op\[2\] as2650.alu_op\[1\] _05772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__11287__A1 _03285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08706_ _02059_ _02976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09686_ _02850_ _03803_ _03847_ _00533_ _03848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_2106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06898_ _01335_ _01338_ _01058_ _01339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_55_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08152__A1 _02327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07561__I _01988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08637_ _01822_ _02909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05849_ _05681_ _05690_ _05695_ _05698_ _05702_ _05703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
XTAP_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08568_ _00923_ _02841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07519_ as2650.stack\[15\]\[13\] _01832_ _01819_ as2650.stack\[12\]\[13\] _01950_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_54_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08499_ _02008_ _02772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_22_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08455__A2 _02726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06466__A1 _00911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10530_ _04642_ _04643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10262__A2 _02606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08392__I _02670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout87 net65 net87 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_195_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_86_wb_clk_i_I clknet_4_2_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10461_ _04559_ _04569_ _04574_ _04332_ _04363_ _04575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_148_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09404__A1 as2650.stack\[6\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06218__A1 _00472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11211__A1 as2650.stack\[13\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10392_ net21 _04494_ _04501_ _04509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_129_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11211__B2 as2650.stack\[15\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06769__A2 _01111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07966__A1 _00503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12131_ net85 net76 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_174_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__12012__CLK clknet_4_2_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07736__I _02155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09707__A2 _03865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11013_ _00722_ _00979_ _05111_ _01130_ _05112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_49_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10722__B1 _01822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_4020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06941__A2 _01380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11278__A1 as2650.stack\[14\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_161_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11278__B2 as2650.stack\[12\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11915_ _00284_ clknet_leaf_73_wb_clk_i as2650.stack\[5\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_61_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10111__B _03727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08694__A2 _02963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11846_ _00006_ clknet_leaf_55_wb_clk_i as2650.cycle\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_57_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11777_ _00160_ clknet_leaf_82_wb_clk_i as2650.stack\[3\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08446__A2 _02717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_186_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06457__A1 _00468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11450__A1 _01449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10728_ _04829_ _04836_ _04837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10659_ _02858_ _04009_ _04769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_139_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_173_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06209__A1 _00651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07406__B1 _01757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07709__A1 _02104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11505__A2 _00751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10072__I _04225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05983__A3 _00441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07870_ _02256_ _02264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_68_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07185__A2 _01622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08382__A1 _02672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06821_ _01262_ _01263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_112_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11269__A1 _05351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09540_ _03702_ _03703_ _03704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_84_wb_clk_i clknet_4_8_0_wb_clk_i clknet_leaf_84_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_06752_ _01166_ _01183_ _01193_ _01194_ _01195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_114_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07381__I _01815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09471_ _00616_ _03638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06683_ _01119_ _01124_ _01126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_37_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09882__A1 _04024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08685__A2 _02955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08422_ _02684_ _02700_ _02701_ _02703_ _00176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_91_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_145_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10492__A2 _04581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_120_wb_clk_i_I clknet_4_2_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08353_ _02644_ _02653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10448__S _05703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07304_ _01739_ _01740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_71_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10244__A2 _04387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08284_ _00506_ _02004_ _02593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_177_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_149_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07235_ _01580_ _01577_ _01574_ _01672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_34_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_166_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09398__B1 _03584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07166_ _00488_ _00922_ _01603_ _00974_ _01604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_106_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_3_wb_clk_i_I clknet_4_1_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10691__B _04799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07948__A1 as2650.stack\[10\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06117_ _00575_ _00576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07097_ _01506_ _01527_ _01535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_160_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07556__I _01983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_191_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06048_ _05675_ _00485_ _00507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_160_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_173_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11078__I _05165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09807_ _00816_ _03961_ _03966_ _03917_ _03967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_115_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07999_ _02200_ _02366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_87_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06923__A2 _01219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10710__I _04363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_189_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09738_ _03150_ _03762_ _00641_ _03899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08387__I _02219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08125__A1 _02381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08676__A2 _01433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09669_ _03779_ _03832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_76_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11700_ _00083_ clknet_leaf_114_wb_clk_i as2650.stack\[10\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09720__B _00731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output17_I net17 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06151__A3 _00585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11631_ _00014_ clknet_leaf_37_wb_clk_i as2650.r123\[1\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_42_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11432__A1 _01013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10235__A2 _04373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11562_ _00850_ _02768_ _02752_ _05607_ _05608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_19_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10513_ _04540_ _04626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_11493_ _05548_ _00402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_156_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09946__I _00682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10444_ _04376_ _04556_ _04557_ _04558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_104_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_178_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11196__B1 _03653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10375_ _04489_ _04493_ _04495_ _00337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_108_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06370__I _00815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12045_ _00414_ clknet_leaf_7_wb_clk_i net49 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_133_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07167__A2 _01604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08364__A1 _02521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10171__A1 _00723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06914__A2 _05752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08297__I _00749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08116__A1 _02456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09864__A1 _03974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08667__A2 _00792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11120__B1 _05157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_178_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11829_ _00212_ clknet_4_7_0_wb_clk_i as2650.r123_2\[1\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08419__A2 _02697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_109_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06545__I _00988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10226__A2 _03650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11423__A1 _02119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09092__A2 _03313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_131_wb_clk_i clknet_4_0_0_wb_clk_i clknet_leaf_131_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_35_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07020_ _05733_ _01459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06850__A1 _01290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_127_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07376__I _01810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06280__I as2650.cycle\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08971_ _01696_ _03074_ _03211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_102_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07922_ as2650.stack\[11\]\[8\] _02178_ _02305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_170_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09591__I _00799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08355__A1 _02513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07853_ _02250_ _02251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_68_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10162__A1 _00782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06366__B1 _00812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06905__A2 _01345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06804_ _01245_ _01246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_112_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07784_ _01112_ _02191_ _02192_ _02195_ _02196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA__08107__A1 _02449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06735_ _01169_ _00434_ _01167_ _01178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_09523_ _00985_ _03685_ _03686_ _03687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_65_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07044__C _00656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09855__A1 _03957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06669__A1 _01102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09454_ _02087_ _02536_ _03621_ _03626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08935__I _03107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06666_ _01109_ _01110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_149_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08405_ _01770_ _02138_ _02692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_52_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09385_ _02272_ _03024_ _03218_ _03576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_06597_ net8 _01041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09607__A1 _00538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10217__A2 _02808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08336_ _02632_ _02640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11414__A1 _03558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08267_ _05698_ _02570_ _02574_ _02575_ _02576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_193_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07218_ _01634_ _01654_ _01655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_165_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06841__A1 _01255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08198_ _02516_ _02508_ _02512_ _02518_ _00137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_134_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07149_ _01341_ _01585_ _01586_ _01573_ _01587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_133_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_84_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07286__I _01717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10160_ _02552_ _00555_ _04311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_160_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10091_ _04242_ _04206_ _04244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_134_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08346__A1 as2650.stack\[3\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10440__I _03665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09006__I _02118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10993_ _05088_ _05090_ _03755_ _05092_ _05093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_95_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08649__A2 _01809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09846__B2 _04004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_128_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_167_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_141_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11614_ _05653_ _05654_ _05655_ _05656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__09074__A2 _03067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07085__A1 _05759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11545_ _02847_ _02770_ _05591_ _05592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_89_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08821__A2 _03067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08580__I _02852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11476_ _00729_ _05532_ _05535_ _05536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__11918__CLK clknet_leaf_72_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10427_ as2650.stack\[1\]\[0\] _01789_ _01793_ as2650.stack\[0\]\[0\] _04541_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_152_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10358_ _03649_ _04476_ _04478_ _04479_ _04480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_83_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10392__A1 net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_174_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10289_ _04422_ _04425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_80_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12028_ _00397_ clknet_leaf_41_wb_clk_i as2650.r123\[2\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_6_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10144__A1 _00673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09837__A1 net34 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06520_ _00862_ _05680_ _00964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_98_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07312__A2 _01740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06451_ _00686_ _00896_ _00897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__11181__I _05124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_194_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09170_ _03390_ _03391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_72_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06275__I _00470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06382_ _00653_ _00828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_109_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08121_ as2650.stack\[0\]\[6\] _02445_ _02460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_175_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_50_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09586__I _00778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08704__B _02718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10953__C _00727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08052_ _02174_ _02392_ _02397_ _02408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_134_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07003_ _01309_ _01284_ _01443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_134_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_192_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10383__A1 net46 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08954_ _01602_ _03192_ _03193_ _03194_ _03195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_88_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08328__A1 as2650.stack\[4\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_116_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07905_ _02280_ _02292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_4619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08885_ _01206_ _03108_ _03130_ as2650.r123_2\[1\]\[1\] _03131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_116_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10686__A2 _05737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_99_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07836_ _02046_ _02241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07767_ _02118_ _02181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_71_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09506_ net25 _03671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_129_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06718_ _01159_ _01160_ _01161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_129_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07698_ _02104_ _02119_ _01997_ _02120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_53_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08500__A1 _02341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06649_ _01090_ _00592_ _01092_ _01093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_25_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09437_ _02533_ _03612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__11091__I _05124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_123_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09368_ as2650.stack\[3\]\[4\] _03546_ _03563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_138_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08319_ _02626_ _02627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_103_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09299_ _03509_ _03502_ _03510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_138_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08803__A2 _02475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06814__A1 _01138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11330_ _05421_ _05422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_120_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06290__A2 _00705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11040__B _05137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11261_ _02724_ _04837_ _05354_ _05355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_84_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_106_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08567__A1 _02811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10212_ _03647_ _00700_ _04361_ _04362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_122_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11192_ _01725_ _04741_ _05286_ _05287_ _05242_ _05288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__10374__A1 net44 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10143_ net92 _04099_ _03728_ _04295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__06042__A2 _00494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07744__I _02148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10074_ _00793_ _04228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10126__A1 net92 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_130_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10677__A2 _04749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05928__I0 as2650.r123\[2\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09531__A3 _02738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08575__I _01271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11626__A1 _05674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10429__A2 _04536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09295__A2 _02673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10976_ _05055_ _04701_ _05075_ _05076_ _00357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_90_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_73_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11740__CLK clknet_leaf_116_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07058__A1 _01485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_178_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06805__A1 _01086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06823__I _05766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06805__B2 _01088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11528_ _04462_ _05575_ _05571_ _05540_ _05576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_89_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10601__A2 _04702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11459_ _05517_ _03491_ _05519_ _00397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_125_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08558__A1 _02819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07230__A1 as2650.holding_reg\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input8_I io_in[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05951_ _05760_ _05727_ _05805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10117__A1 _03721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08670_ _02065_ _02848_ _01435_ _02089_ _02942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05882_ _05712_ _05736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__09522__A3 _00986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10668__A2 _01738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07533__A2 _01961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07621_ _01984_ _01998_ _02026_ _02048_ _00030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_26_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07552_ _01980_ _01728_ _01849_ _01981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__10948__C _00673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11617__A1 _05638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06503_ _00945_ _00946_ _00947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07483_ as2650.stack\[5\]\[12\] _01914_ _01856_ as2650.stack\[4\]\[12\] _01915_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_107_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09222_ _03436_ _03440_ _03441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_139_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05847__A2 _05693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06434_ _00879_ _00880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_33_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09153_ as2650.r123_2\[2\]\[1\] _03342_ _03374_ _03163_ _03375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_104_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06365_ _00550_ _00713_ _00721_ _00812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_104_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08104_ _02394_ _02436_ _02444_ _02447_ _00114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08797__A1 _03044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07829__I net71 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09084_ _01641_ _01653_ _03307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_148_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06296_ _00485_ _00748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_190_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_147_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08035_ _02050_ _02394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06272__A2 _00717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08549__A1 _02345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_150_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10356__A1 _00881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06024__A2 _00482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09986_ _04137_ _04141_ _04142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_5117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07564__I net73 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07772__A2 _02178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08937_ _02836_ _03080_ _03179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_150_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11305__B1 _05303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11086__I _00755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10659__A2 _04009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08868_ _03081_ _03114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08721__A1 _02405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08721__B2 _02987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07819_ _02226_ _02227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_2_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06732__B1 _01173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11961__D _00330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08799_ as2650.stack\[8\]\[6\] _03026_ _03048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10830_ _02619_ _04921_ _04935_ _04936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__11608__A1 _02778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08395__I _02230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09277__A2 _03491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11763__CLK clknet_leaf_80_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10761_ _04237_ _04866_ _04868_ _04869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_183_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10692_ _02105_ _03957_ _02080_ _04653_ _04801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_8_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_157_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_194_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08788__A1 _03037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10595__A1 _04596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08252__A3 _00873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_193_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07460__A1 _01854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11313_ as2650.stack\[13\]\[6\] _05171_ _05310_ as2650.stack\[15\]\[6\] _05406_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_154_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11244_ as2650.stack\[14\]\[4\] _05180_ _05269_ as2650.stack\[12\]\[4\] _05215_ _05339_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_106_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05861__I2 as2650.r123_2\[1\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09201__A2 _01517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11544__B1 _04429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07063__I1 _01501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11175_ as2650.stack\[9\]\[2\] _05266_ _05272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08960__A1 _01619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10126_ net92 _04277_ _04278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_136_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_23_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10057_ _04209_ _04210_ _04211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_5684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09903__B _03968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08712__A1 as2650.stack\[15\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_149_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09268__A2 _03338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07279__A1 _00947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10959_ _02229_ _00628_ _00779_ _05060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_189_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08779__A1 _03028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_38_wb_clk_i clknet_4_6_0_wb_clk_i clknet_leaf_38_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_145_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06150_ _00489_ _00594_ _00609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_160_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_185_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10586__A1 _04620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07451__A1 _01263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06081_ _00531_ _00540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06254__A2 _00697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_172_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_37_wb_clk_i_I clknet_4_6_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_173_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11636__CLK clknet_leaf_39_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07203__A1 _05723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06006__A2 _00462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09840_ _02105_ _01464_ _03999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_98_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07384__I _01818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09771_ _00728_ _03931_ _00297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06983_ _00430_ _05808_ _00434_ _05770_ _01423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_140_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_189_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08722_ as2650.stack\[15\]\[5\] _02978_ _02988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09813__B _03972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05934_ as2650.ins_reg\[4\] as2650.alu_op\[0\] _05788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_6_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11786__CLK clknet_leaf_85_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_167_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05865_ _05718_ _05719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_96_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08653_ _02805_ _02924_ _02776_ _02925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_54_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10510__A1 as2650.stack\[7\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10510__B2 as2650.stack\[5\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10678__C _04744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07604_ _05675_ _02018_ _02032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_148_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08584_ _02845_ _02847_ _02851_ _02856_ _02857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_148_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07535_ as2650.stack\[3\]\[14\] _01912_ _01856_ as2650.stack\[0\]\[14\] _01859_ as2650.stack\[1\]\[14\]
+ _01965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_169_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10813__A2 _04915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07466_ as2650.stack\[15\]\[11\] _01874_ _01877_ as2650.stack\[14\]\[11\] _01899_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_74_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06664__S _05710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10694__B _02107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09205_ _03414_ _03424_ _03425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06417_ _00862_ _00863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_leaf_76_wb_clk_i_I clknet_4_11_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07397_ _01810_ _01832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_176_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09136_ _01646_ _03357_ _03358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_148_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06348_ _00777_ _00797_ _00008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10577__A1 as2650.stack\[9\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10577__B2 as2650.stack\[8\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09067_ _03202_ _03257_ _03291_ _03292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_120_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06279_ _00707_ _00732_ _00733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_151_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_163_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07993__A2 _02360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08018_ _02181_ _02202_ _02356_ _02380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_150_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09707__C _03728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09195__A1 _05759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09734__A3 _01285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06412__B _00609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08942__A1 _01954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11541__A3 _05571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09969_ _04075_ _01695_ _04125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_4202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_134_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09498__A2 _03660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_output47_I net47 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11931_ _00300_ clknet_leaf_62_wb_clk_i net36 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_4279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_57_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_175_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08170__A2 _02497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10588__C _04645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07243__B _00825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11862_ _00231_ clknet_leaf_27_wb_clk_i as2650.r123_2\[0\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06638__I _01081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10813_ _04654_ _04915_ _04918_ _04651_ _04919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_26_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11793_ _00176_ clknet_leaf_86_wb_clk_i as2650.stack\[1\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10744_ _00894_ _04851_ _04852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__10804__A2 _04470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10675_ _04780_ _04781_ _04784_ _04785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_40_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11212__C _05215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10568__A1 _00517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06236__A2 _00580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07433__A1 as2650.stack\[2\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_142_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07984__A2 _02352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_181_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09186__B2 _03163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11227_ _02927_ _05130_ _00847_ _05322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_136_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08933__A1 _03110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06539__A3 _00982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11158_ _00426_ _00680_ _03782_ _05240_ _05254_ _05255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__10740__A1 _04229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10109_ _04249_ _04261_ _04262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_11089_ _01102_ _05125_ _05187_ _05188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_5470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09489__A2 _01712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06548__I _00743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06172__A1 _00536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08700__A4 _02023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07320_ _01755_ _01756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_147_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_147_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07251_ _01600_ _01687_ _01688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_143_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07672__A1 _02094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_158_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06202_ _00647_ _00660_ _00661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_14_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07182_ _01288_ _01619_ _01620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__06283__I _00736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_191_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10559__A1 _03790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09413__A2 _02514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06133_ _00591_ _00592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06227__A2 _05680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10023__A3 _04120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07975__A2 net77 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06064_ _00456_ _00523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09177__A1 _05732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08924__A1 _03165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09823_ _01466_ _01458_ _03981_ _03982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_134_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10326__A4 _04340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11523__A3 _05571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09754_ _00881_ _00730_ _03915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06966_ _01402_ _01335_ _01404_ _01405_ _01406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_39_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10689__B _04586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08705_ _02384_ _02970_ _02973_ _02975_ _00187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05917_ as2650.alu_op\[0\] _05771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11287__A2 _05189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09685_ _03842_ _03845_ _03846_ _03847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_54_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06897_ _01237_ _01239_ _01245_ _01338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_54_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08152__A2 _02480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08636_ _02781_ _02908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05848_ _05700_ _05701_ _05702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07360__B1 _01795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_120_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08567_ _02811_ _02832_ _02839_ _02840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_184_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09101__A1 _05764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07518_ as2650.stack\[14\]\[13\] _01812_ _01816_ as2650.stack\[13\]\[13\] _01949_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_19_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10798__A1 _04610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08498_ _02747_ _02337_ _02769_ _02770_ _02771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_161_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08455__A3 _02727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout88 net64 net88 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07449_ _01777_ _01883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_183_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10460_ _03723_ _04570_ _04573_ _04574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_167_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09404__A2 _03585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09119_ _03098_ _03298_ _03341_ _00235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_135_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06218__A2 _00673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10391_ _03285_ _04490_ _04507_ _04508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_136_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11211__A2 _05266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08622__B _02894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12130_ net81 net14 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_159_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07966__A2 _01087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11951__CLK clknet_leaf_49_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05977__A1 _00428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10970__A1 _03749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09168__A1 _05723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_152_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08915__A1 _01303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11012_ _00533_ _00973_ _00986_ _05111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_81_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10722__A1 as2650.stack\[11\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10722__B2 as2650.stack\[10\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_77_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_161_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11278__A2 _01933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_161_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08143__A2 _02477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09340__A1 as2650.stack\[4\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11914_ _00283_ clknet_leaf_73_wb_clk_i as2650.stack\[5\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_18_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11845_ _00005_ clknet_leaf_54_wb_clk_i as2650.cycle\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_45_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09900__C _03917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08583__I _02855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11776_ _00159_ clknet_leaf_82_wb_clk_i as2650.stack\[3\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_14_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10789__A1 _02902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06457__A2 _00550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07654__A1 as2650.stack\[13\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10727_ _01844_ _04832_ _04835_ _04836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__11450__A2 _05499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_186_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10658_ _03960_ _04767_ _04768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_127_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06209__A2 _00667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07406__A1 as2650.stack\[14\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07406__B2 as2650.stack\[12\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10589_ _04642_ _04700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_142_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07957__A2 _02278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10961__A1 _00784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07148__B _01346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07709__A2 _02129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08382__A2 _02667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06820_ _01210_ _01262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_110_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06393__A1 _00590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07662__I _02086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06751_ _01166_ _01178_ _01194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09331__A1 as2650.stack\[4\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_184_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06682_ _01119_ _01124_ _01125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_09470_ _00899_ _00758_ _03637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_64_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06278__I _00731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08685__A3 _02956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08421_ as2650.stack\[1\]\[13\] _02697_ _02703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_36_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07893__A1 as2650.stack\[10\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09810__C _03883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11824__CLK clknet_leaf_100_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_53_wb_clk_i clknet_4_13_0_wb_clk_i clknet_leaf_53_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_08352_ _02505_ _02646_ _02647_ _02652_ _00157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_177_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05910__I as2650.r0\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07303_ _01738_ _01739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08283_ _00649_ _02592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_32_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07234_ _01669_ _01670_ _01671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_14_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11974__CLK clknet_leaf_49_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09398__A1 _03555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07165_ _00928_ _00558_ _01603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_118_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_145_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06116_ _00535_ _00561_ _00575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07948__A2 _02319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08070__A1 _02153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07096_ _01506_ _01527_ _01534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_145_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_156_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10952__A1 as2650.ivec\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10952__B2 _05028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06047_ _00505_ _00506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_132_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10704__A1 _04808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09806_ _03951_ _03867_ _03965_ _03966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_25_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07998_ _02187_ _02365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07572__I _01993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09737_ _02854_ _01322_ _03897_ _03898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__11308__B _05265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06949_ _01237_ _01239_ _01342_ _01333_ _01245_ _01389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_55_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09322__A1 as2650.stack\[4\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06188__I _00542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09668_ _03787_ _03815_ _03829_ _03830_ _03831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__06136__A1 _00589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_182_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08619_ _02778_ _02804_ _02871_ _02891_ _02892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XTAP_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07884__A1 as2650.stack\[10\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09599_ _03762_ _03763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09499__I _00929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10866__C _04298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11630_ _05665_ _05667_ _05668_ _00712_ _00419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__07521__B _01951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05820__I _05673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11432__A2 _00934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10235__A3 _04383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11561_ _00863_ _02732_ _00613_ _05131_ _05607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_156_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_180_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10512_ _02907_ _04623_ _04624_ _04625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_155_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11492_ as2650.r123\[3\]\[3\] _05548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_149_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_155_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09389__A1 _02045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10443_ _03722_ _00779_ _04557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_6_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09448__B _03621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11196__A1 _01269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_193_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11196__B2 _02856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08061__A1 _02412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10374_ net44 _04494_ _04301_ _04495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_136_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10943__A1 _04242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06611__A2 _00987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12044_ _00413_ clknet_4_4_0_wb_clk_i net52 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_172_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_78_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_117_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08578__I _02850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06375__A1 _00472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10171__A2 _04308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06375__B2 _00446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07482__I _01830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08116__A2 _02425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09313__A1 _02388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06098__I _00466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_185_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11120__A1 as2650.stack\[2\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11120__B2 as2650.stack\[0\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07875__A1 as2650.stack\[12\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05886__B1 _05738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11828_ _00211_ clknet_leaf_34_wb_clk_i as2650.r123_2\[1\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_159_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10226__A3 _01131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11759_ _00142_ clknet_leaf_82_wb_clk_i as2650.stack\[5\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_18_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11423__A2 _05462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06850__A2 _01291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11187__A1 _05238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07657__I _02081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08052__A1 _02174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_170_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10934__A1 _04395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10083__I _00800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08970_ _02345_ _03111_ _03209_ _03210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_130_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_100_wb_clk_i clknet_4_3_0_wb_clk_i clknet_leaf_100_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_102_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05956__A4 _05769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07921_ _02160_ _02304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_29_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07852_ _01985_ _02031_ _02249_ _02250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_60_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06366__A1 _00811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06366__B2 _00639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10162__A2 _02737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07392__I _01826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05905__I _05758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06803_ _01233_ _01245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput1 io_in[10] net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_84_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07783_ _02194_ _02195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_37_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09304__A1 _03044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09522_ _01005_ _00905_ _00986_ _03686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_06734_ _00885_ _01176_ _01177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__06118__A1 _00523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09855__A2 _01435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07866__A1 _02214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09453_ as2650.stack\[5\]\[3\] _03615_ _03625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06665_ _01108_ _01109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_1854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08404_ as2650.stack\[1\]\[8\] _02689_ _02691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_149_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12002__CLK clknet_4_15_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09384_ _03574_ _03575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09607__A2 _00723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06596_ _01039_ _01040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_40_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08335_ _02627_ _02639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_71_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07060__C _01166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10217__A3 _00496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11414__A2 _05473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09083__A3 _01652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08951__I _03115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08266_ _00886_ _00686_ _02575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08291__A1 _00506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07217_ _01641_ _01653_ _01654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_137_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06841__A2 _01256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08197_ as2650.stack\[6\]\[10\] _02517_ _02518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__11178__A1 _05271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08043__A1 _02167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07148_ _01082_ _01585_ _01346_ _01586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11310__C _05174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07079_ _01517_ _01518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_161_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10090_ _04242_ _04203_ _04243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_121_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09543__A1 _00747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08346__A2 _02645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08398__I _02236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11350__A1 _05222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05815__I as2650.cycle\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09731__B _00533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10992_ _04439_ _05084_ _05091_ _04364_ _05092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_16_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07857__A1 _02154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_188_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10596__C _04604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06646__I _05695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_160_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11613_ _05638_ _04440_ _04441_ _05185_ _05655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_184_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08861__I _03107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08282__A1 _00852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11544_ _05672_ _00861_ _05589_ _04429_ _05522_ _05591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_89_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_123_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11475_ _04524_ _05534_ _05535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_7_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07477__I as2650.r123\[0\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06381__I _05693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08034__A1 _02384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10426_ _02788_ _04540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_125_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08034__B2 _02393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10916__A1 _04610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09782__A1 _02859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10357_ _04326_ _03637_ _04380_ _03659_ _04479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_112_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10288_ _04424_ _00321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08337__A2 _02636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09534__A1 _03687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12027_ _00396_ clknet_leaf_39_wb_clk_i as2650.r123\[2\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_26_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10631__I _02758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11341__A1 _05216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05946__I1 _05786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__12025__CLK clknet_leaf_39_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07848__A1 _02053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_165_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06556__I _00968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06450_ _00895_ _00896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_61_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_181_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06520__A1 _00862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06381_ _05693_ _00827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_37_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09867__I _02826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08120_ _02409_ _02454_ _02458_ _02459_ _00118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_147_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10080__A1 _04209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08051_ as2650.stack\[12\]\[4\] _02390_ _02407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07387__I _01779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07002_ _01430_ _01264_ _01013_ _01441_ _01442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__06291__I as2650.cycle\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10907__A1 _04596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06587__A1 net50 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11580__A1 _01327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08953_ _01611_ _03114_ _03192_ _03194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_9_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09525__A1 _00772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08328__A2 _02634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07904_ _02078_ _02270_ _02290_ _02291_ _00070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_69_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08884_ _03104_ _03130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_29_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07835_ as2650.stack\[13\]\[8\] _02104_ _02240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_3919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07766_ as2650.stack\[11\]\[6\] _02163_ _02180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09043__S _03271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09505_ _01091_ _03669_ _03670_ _00292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_53_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06717_ _01119_ _01158_ _01160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__07839__A1 as2650.stack\[13\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07697_ _02118_ _02119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_64_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_169_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08500__A2 _02566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09436_ _01980_ _03601_ _03611_ _00282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06648_ _01080_ _01091_ _01092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09367_ _02651_ _03562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06579_ _01022_ _00944_ _01023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_166_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11399__A1 _02003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08318_ _01985_ _02485_ _02486_ _02626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__07067__A2 _01382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08264__A1 _00686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09298_ _02096_ _03509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_90_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_193_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06814__A2 _00432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08249_ _02557_ _02558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_193_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_165_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08016__A1 _02102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11040__C _05138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11260_ _05352_ _05353_ _02814_ _00842_ _05354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_137_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10211_ _04331_ _00786_ _04103_ _04361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_106_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11191_ _02000_ _00874_ _05192_ _05287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_121_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11571__A1 _02956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output77_I net77 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10142_ _00810_ _04293_ _04294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09516__A1 _00648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10073_ _04223_ _03752_ _04224_ _04226_ _04227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_153_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11323__A1 _04409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12048__CLK clknet_leaf_9_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08856__I _03102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09461__B _03612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06750__A1 _01188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06750__B2 _01058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11626__A2 _04394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10975_ _04404_ _05076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_189_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_44_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06376__I _00731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_160_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09687__I _00980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08255__A1 _02561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10062__A1 net66 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11231__B _05325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11527_ _05570_ _05575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_195_1819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08007__A1 _02170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_27_wb_clk_i_I clknet_4_7_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11458_ _01707_ _05502_ _05513_ as2650.r123\[2\]\[7\] _05519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_171_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10409_ _02732_ _00705_ _04521_ _04522_ _04523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_139_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_3_4_0_wb_clk_i clknet_0_wb_clk_i clknet_3_4_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_67_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06569__A1 _01001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11389_ _05460_ _05468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_152_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11562__A1 _00850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_139_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_171_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09507__A1 _00483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10361__I _04482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05950_ _05802_ _05803_ _05804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_112_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07518__B1 _01816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11314__A1 _05177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05881_ _05733_ _05734_ _05735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07620_ _02036_ _02045_ _02047_ _02048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08730__A2 _02978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07670__I _02093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07551_ _01664_ _01980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_35_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11617__A2 _04429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06502_ _00924_ _00946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_35_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06286__I _00711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07482_ _01830_ _01914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_50_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08494__A1 _02752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09221_ _01569_ _02233_ _03440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06433_ _00878_ _00879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_72_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_66_wb_clk_i_I clknet_4_12_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09152_ _03344_ _03373_ _03374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_147_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06364_ _00810_ _00811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_175_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10053__A1 _04200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08103_ as2650.stack\[0\]\[1\] _02445_ _02446_ _02447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_147_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08797__A2 _03041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09083_ _01547_ _01551_ _01652_ _03306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_147_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06295_ _00746_ _00747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_120_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_159_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08034_ _02384_ _02386_ _02391_ _02393_ _00098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_176_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09746__A1 _02081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08549__A2 _02821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_192_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10356__A2 _00611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11553__A1 _05108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09985_ _04047_ _04139_ _04140_ _04141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_115_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08936_ _03096_ _03178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_103_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_4406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11305__A1 as2650.stack\[0\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06980__A1 _01390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11305__B2 as2650.stack\[3\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08867_ _03079_ _03113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08721__A2 _02985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07818_ _02223_ _02190_ _02124_ _02225_ _02226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_85_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08798_ _02112_ _03047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_44_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11069__B1 _05163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11608__A2 _04786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07749_ _02073_ _02167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_77_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_26_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08485__A1 _00798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10760_ _03642_ _04859_ _04867_ _04819_ _04868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_148_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09419_ as2650.ivec\[0\] _01102_ _03601_ _03602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_125_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10691_ _04794_ _04793_ _04799_ _04800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_70_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08237__A1 _00898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08788__A2 _03022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_165_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_154_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06145__B _00509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10595__A2 _04704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08252__A4 _02555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11312_ as2650.stack\[14\]\[6\] _05268_ _01961_ as2650.stack\[12\]\[6\] _05405_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_148_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_153_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09737__A1 _02854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11243_ as2650.stack\[13\]\[4\] _05266_ _05172_ as2650.stack\[15\]\[4\] _05338_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_88_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05861__I3 as2650.r123_2\[0\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08360__B _02652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11544__A1 _05672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11174_ _05267_ _05270_ _05271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10125_ _04256_ _04246_ _04277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10181__I _04331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06971__A1 _01077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10056_ net39 net38 _04133_ _04210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_5674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_102_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08712__A2 _02972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08586__I _02858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_100_wb_clk_i_I clknet_4_3_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07279__A2 _00953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08476__A1 _02745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10958_ _04814_ _05046_ _05057_ _04794_ _05059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_182_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10283__A1 _00941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10889_ _04879_ _04985_ _04990_ _04771_ _04992_ _04993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_73_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08228__A1 _02519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10035__A1 _04181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_129_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08779__A2 _03022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_184_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10586__A2 _04649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06080_ _00529_ _00534_ _00538_ _00539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__06254__A3 _00708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11535__A1 _04462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07203__A2 _01109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06006__A3 _00464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08400__A1 _02686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09770_ _03886_ _03837_ _03930_ _03931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_101_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06982_ _01421_ _01422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06962__A1 _01230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08721_ _02405_ _02985_ _02986_ _02987_ _00191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__11299__B1 _05390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05933_ as2650.alu_op\[2\] _05692_ _05787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09900__A1 _00810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08652_ _02912_ _02917_ _02923_ _01845_ _02924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_67_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05864_ _05717_ _05718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_94_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10510__A2 _01835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07603_ _01994_ _02031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08583_ _02855_ _02856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_78_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06190__A2 _00593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07534_ _01854_ _01960_ _01963_ _01964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_81_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10274__A1 _00978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07465_ as2650.stack\[11\]\[11\] _01858_ _01872_ _01898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_179_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09204_ _03389_ _03423_ _03424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_33_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06416_ as2650.prefixed _00862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_195_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07396_ as2650.stack\[2\]\[9\] _01824_ _01827_ as2650.stack\[0\]\[9\] _01830_ as2650.stack\[1\]\[9\]
+ _01831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_52_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09135_ _05750_ _01649_ _03357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_147_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06347_ _00611_ _00644_ _00796_ _00797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_124_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_159_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10577__A2 _01790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09066_ _01974_ _03251_ _03278_ _03290_ _03291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_06278_ _00731_ _00732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08017_ as2650.stack\[14\]\[6\] _02362_ _02379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_135_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_151_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07575__I _02002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10215__B _04364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08942__A2 _03111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09968_ _04034_ _04037_ _04123_ _04082_ _04124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_76_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_89_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08919_ _03103_ _03163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_4214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09899_ _04041_ _03820_ _04057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_111_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10869__C _04912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11930_ _00299_ clknet_leaf_62_wb_clk_i net35 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_4258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06705__A1 _01146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10501__A2 _04612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05823__I _05676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11861_ _00230_ clknet_leaf_30_wb_clk_i as2650.r123_2\[0\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_168_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_26_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10812_ _04916_ _04917_ _04918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08458__A1 _02730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11792_ _00175_ clknet_leaf_86_wb_clk_i as2650.stack\[1\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10885__B _04897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10743_ _04849_ _04797_ _04847_ _04848_ _04851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_9_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08355__B _02652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_186_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10674_ _01732_ _04782_ _04783_ _04784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_139_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09958__A1 _04087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_185_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10176__I _04326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06236__A3 _00684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07433__A2 _01865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09186__A2 _03342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11226_ _05200_ _01422_ _05319_ _05320_ _03859_ _05321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_136_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09430__I0 as2650.ivec\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08933__A2 _03174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11157_ _02841_ _03815_ _05252_ _05253_ _05254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_81_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10740__A2 _05746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10108_ _04250_ _04260_ _04261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11088_ _05147_ _05148_ _05186_ _05187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_5471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10039_ _04109_ _04189_ _04190_ _04193_ _04194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__07434__B _01846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06829__I net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08697__A1 _02905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_149_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_125_wb_clk_i clknet_4_0_0_wb_clk_i clknet_leaf_125_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__06172__A2 as2650.cycle\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11453__B1 _05513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10287__S _04423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07121__A1 _01541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07250_ _05797_ _01454_ _01687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_56_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10008__A1 _02195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06201_ _00648_ _00650_ _00659_ _00660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_31_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09949__A1 _03866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11205__B1 _05297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07181_ _01618_ _01619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09949__B2 _04087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_185_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10559__A2 _05782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_195_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06132_ _00453_ _05692_ _00591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_145_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06063_ _00521_ _00522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07395__I _01829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09177__A2 _01517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11753__CLK clknet_leaf_81_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09421__I0 as2650.ivec\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09822_ _03937_ _03979_ _03938_ _03980_ _03981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_141_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10731__A2 _04793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_189_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09753_ _02080_ _03914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06965_ _01342_ _01326_ _01405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_171_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08704_ _02276_ _02974_ _02718_ _02975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05916_ _05769_ _05770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09684_ _03842_ _03845_ _01002_ _03846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_27_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06896_ _01335_ _01336_ _01337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_3_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08635_ _02906_ _02907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05847_ _05691_ _05693_ _05701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_55_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07360__B2 as2650.stack\[12\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08566_ _02833_ _01700_ _02838_ _02839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_23_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10247__A1 _04391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09101__A2 _01515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07517_ as2650.stack\[10\]\[13\] _01944_ _01866_ _01948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_195_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07112__A1 _05765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08497_ _02348_ _02615_ _02770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_74_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11380__I _05455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08455__A4 _00883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07448_ _01871_ _01873_ _01881_ _01882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__06466__A3 _00703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07663__A2 _02087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout89 net57 net89 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_10_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07379_ _01750_ _01814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_148_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09118_ _03108_ _03337_ _03340_ as2650.r123_2\[2\]\[0\] _03341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_148_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07415__A2 _01847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10390_ _02835_ _04491_ _04507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09049_ _03276_ as2650.r123_2\[0\]\[3\] _03271_ _03277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_139_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05818__I _05671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09168__A2 _01380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_26_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11011_ _00941_ _02759_ _00637_ _05110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_117_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10722__A2 _04822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10486__A1 _04597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11913_ _00282_ clknet_leaf_69_wb_clk_i as2650.ivec\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_79_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11844_ _00000_ clknet_leaf_67_wb_clk_i as2650.cycle\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11775_ _00158_ clknet_leaf_92_wb_clk_i as2650.stack\[3\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_53_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07103__A1 _05776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10789__A2 _04889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08085__B _02431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06384__I _00829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10726_ _02906_ _04833_ _04834_ _04835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__06457__A3 _00713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07654__A2 _02025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10657_ _04764_ _04765_ _04763_ _04721_ _04767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__08813__B _03057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11776__CLK clknet_leaf_82_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07406__A2 _01781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10588_ _02071_ _04531_ _04699_ _04645_ _00346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_157_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10410__A1 _00662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10961__A2 _00681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11209_ _05216_ _05301_ _05304_ _05305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_110_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07943__I _02206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_68_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06393__A2 _05695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07590__A1 _02004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06750_ _01188_ _01190_ _01192_ _01058_ _01193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_49_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09331__A2 _03521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06681_ _01120_ _01122_ _01123_ _01124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_97_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06145__A2 _00603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08420_ _02680_ _02700_ _02701_ _02702_ _00175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_64_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08774__I _02050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07893__A2 _02274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08351_ _02651_ _02652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_166_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07302_ _01737_ _01738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06294__I as2650.cycle\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08282_ _00852_ _00861_ _02591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08842__A1 _01100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07233_ _01662_ _01668_ _01670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_105_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_93_wb_clk_i clknet_4_8_0_wb_clk_i clknet_leaf_93_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_30_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_30_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09398__A2 _03575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07164_ _01601_ _01602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06115_ _00524_ _00574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_173_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07095_ _01504_ _01529_ _01532_ _01533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_105_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08070__A2 _01989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06046_ _00487_ _00504_ _00505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_133_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06908__A1 _01327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10704__A2 _04810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07853__I _02250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09805_ _00629_ _03964_ _03965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_64_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07997_ _02059_ _02364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_75_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07581__A1 _00518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07581__B2 _02008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06948_ as2650.r123\[1\]\[4\] _01116_ _01387_ _01223_ _01388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_09736_ _03851_ _03895_ _03896_ _03897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_101_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_186_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09667_ _00451_ _03830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_27_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06879_ _01269_ _01284_ _01320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_131_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11649__CLK clknet_leaf_134_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06136__A2 _05787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08618_ _02885_ _02888_ _02890_ _02891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08684__I _02597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09598_ _01128_ _03762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_27_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07884__A2 _02274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_184_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08549_ _02345_ _02821_ _02590_ _02822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11799__CLK clknet_leaf_121_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11560_ _05599_ _05604_ _05605_ _05606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__11432__A3 _01055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_128_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10511_ as2650.stack\[6\]\[1\] _01823_ _01794_ as2650.stack\[4\]\[1\] _04624_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_126_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10640__A1 _02093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11491_ _05547_ _00401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_137_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08633__B _00647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10442_ _04076_ _03731_ _04555_ _04556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09389__A2 _03579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11196__A2 _02866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08352__C _02652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10373_ _04480_ _04494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_48_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08061__A2 _02406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06611__A3 _00995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_151_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12043_ _00412_ clknet_4_4_0_wb_clk_i net78 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09464__B _03612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09010__A1 _02302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07763__I _02155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06914__A4 _01212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06379__I _00491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07324__A1 _01735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11120__A2 _05212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08594__I _02866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05886__B2 _05739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11827_ _00210_ clknet_leaf_106_wb_clk_i as2650.stack\[8\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11758_ _00141_ clknet_leaf_80_wb_clk_i as2650.stack\[6\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_124_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10709_ _02351_ _04792_ _04818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11689_ _00072_ clknet_leaf_0_wb_clk_i as2650.stack\[10\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07938__I _02196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_155_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_161_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11187__A2 _03147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08052__A2 _02392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10934__A2 _03824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_142_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06998__B _01035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07920_ _02122_ _02292_ _02301_ _02303_ _00074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_69_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09001__A1 _03040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_116_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08769__I _02022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11344__C1 as2650.stack\[10\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07673__I _02096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_190_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07851_ _02033_ _02249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09552__A2 _02584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06366__A2 _00717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06802_ _01242_ _01243_ _01244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_112_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10162__A3 _03678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_68_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput2 io_in[11] net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07782_ _02193_ _02194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10032__C _04105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09521_ _02552_ _00547_ _03685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_83_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06733_ as2650.holding_reg\[1\] _01168_ _01173_ _01176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__09304__A2 _03508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06118__A2 _00574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10967__C _02350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09452_ _03555_ _03613_ _03623_ _03624_ _00285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06664_ as2650.r123\[0\]\[0\] as2650.r123_2\[0\]\[0\] _05710_ _01108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_1844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06669__A3 _01112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07866__A2 _02252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__11941__CLK clknet_leaf_56_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08403_ _02689_ _02690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_40_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09068__A1 as2650.r123_2\[0\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10870__A1 net65 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10539__I _02350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09383_ _02510_ _03574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_51_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06595_ _00947_ _01038_ _01039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_40_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08334_ _02519_ _02628_ _02633_ _02638_ _00153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_127_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08009__I _02200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10217__A4 _00787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_178_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10622__A1 as2650.stack\[3\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08265_ _05670_ _00735_ _02574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_119_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08291__A2 _02599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07216_ _01642_ _01652_ _01653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_20_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08196_ _02506_ _02517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_152_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07147_ _01574_ _01585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_101_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08043__A2 _02392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_156_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07078_ _01516_ _01517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_66_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_153_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06029_ _00487_ _00448_ _00488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_133_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08679__I net54 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09543__A2 _00546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09719_ _03874_ _03875_ _03880_ _03881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_56_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10991_ _03816_ _05080_ _05091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_27_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10877__C _04891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_4_6_0_wb_clk_i clknet_3_3_0_wb_clk_i clknet_4_6_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07857__A2 _02136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output22_I net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05831__I _05684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05868__A1 _05720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10861__A1 _04752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11612_ _02805_ _04741_ _05654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_168_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_141_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10613__A1 _02855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_180_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11543_ _05156_ _05162_ _05590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_129_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08282__A2 _00861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07758__I _02096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06662__I _01105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11474_ _00740_ _02599_ _05533_ _00519_ _05534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__07490__B1 _01879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_184_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_clkbuf_leaf_17_wb_clk_i_I clknet_4_5_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10425_ _01786_ _04537_ _04538_ _04539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_67_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09973__I _03948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10916__A2 _05007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09782__A2 _03803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10356_ _00881_ _00611_ _04477_ _04478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_140_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_139_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11814__CLK clknet_leaf_108_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10287_ _04417_ _01061_ _04423_ _04424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_78_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12026_ _00395_ clknet_leaf_39_wb_clk_i as2650.r123\[2\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_191_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09922__B _03769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07848__A2 _02231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10359__I _04480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06520__A2 _05680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_56_wb_clk_i_I clknet_4_15_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06380_ _00477_ _00826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_1590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_147_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10604__A1 _03150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09470__A1 _00899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07668__I _02046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06284__A1 _00468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08050_ _02256_ _02406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06572__I as2650.addr_buff\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10080__A2 _02955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06284__B2 _00737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07481__B1 _01855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07001_ _01431_ _01307_ _01440_ _01052_ _01441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_116_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09883__I net36 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06036__A1 _00491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06587__A2 _01030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07784__A1 _01112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11580__A2 _01416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07784__B2 _02195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08952_ _05801_ _03059_ _03193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08499__I _02008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05916__I _05769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout89_I net57 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09525__A2 _00784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07903_ _02170_ _02285_ _02286_ _02291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08883_ _03069_ _03126_ _03128_ _03129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_130_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07536__A1 as2650.stack\[2\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07834_ _02052_ _02239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_29_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_170_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_95_wb_clk_i_I clknet_4_9_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07765_ _02102_ _02172_ _02176_ _02179_ _00043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_186_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08448__B _02718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06716_ _01119_ _01158_ _01159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_09504_ net24 _03669_ _02894_ _03670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11096__A1 _01725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07839__A2 _02242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07696_ _02116_ _02083_ _02117_ _02118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_164_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09435_ as2650.ivec\[7\] _03601_ _03611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06647_ _05694_ _01091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08500__A3 _02772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_94_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_36_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09366_ _02090_ _03561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06578_ _01021_ _01022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_36_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11399__A2 _02146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08317_ _02605_ _02623_ _02624_ _02625_ _00149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_193_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08264__A2 _02572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09297_ _02670_ _03508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09461__A1 _02110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08248_ _00470_ _00569_ _02557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_138_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_107_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_180_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09213__A1 _03162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08016__A2 _02373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08179_ _02327_ _02500_ _02501_ _02503_ _00133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
Xclkbuf_opt_1_0_wb_clk_i clknet_4_1_0_wb_clk_i clknet_opt_1_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_118_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10210_ net91 _00971_ _03649_ _04360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__06027__A1 _00483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11020__A1 _03646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11190_ _01028_ _05245_ _05286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_136_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07775__A1 _02186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10141_ _04284_ _04292_ _04293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__10732__I _02557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09516__A2 _02593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11987__CLK clknet_leaf_77_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10072_ _04225_ _04226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08202__I _02226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07246__C _01165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11323__A2 _01693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10531__B1 _04619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_29_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08358__B _02652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11087__A1 _05152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06657__I _01100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10974_ _04532_ _05058_ _05074_ _03757_ _04744_ _05075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_43_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_16_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10834__A1 _04161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_169_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_31_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09452__A1 _03555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08255__A2 _02563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06266__A1 _00531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11231__C _02960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11526_ _05574_ _00409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11457_ _05517_ _03484_ _05518_ _00396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08007__A2 _02202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11011__A1 _00941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10408_ _00602_ _02573_ _04522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08558__A3 _02830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11388_ _05456_ _05467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_152_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06569__A2 _00981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07766__A1 as2650.stack\[11\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11562__A2 _02768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10339_ _04377_ _00887_ _04465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10642__I _02824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_140_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09507__A2 _02554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_87_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07518__A1 as2650.stack\[14\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12009_ _00378_ clknet_leaf_117_wb_clk_i as2650.stack\[9\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_39_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05880_ _05726_ _05734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_39_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10522__B1 _01826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10798__B _04903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11473__I _04525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07550_ as2650.r123\[0\]\[7\] _01979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__06567__I _01010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06501_ _00744_ _00937_ _00945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_59_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_165_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10825__A1 _04116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07481_ as2650.stack\[7\]\[12\] _01912_ _01855_ as2650.stack\[6\]\[12\] _01913_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__09691__A1 _01274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09220_ _03437_ _03438_ _03439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_34_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06432_ _05704_ _00878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_194_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_166_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09151_ _03346_ _03372_ _03373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06363_ _00809_ _00810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09443__A1 _02045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08102_ _02423_ _02446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09082_ _01639_ _01640_ _03304_ _03305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_108_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06294_ as2650.cycle\[8\] _00746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_148_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10038__B _03727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_194_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08033_ _02276_ _02392_ _02264_ _02393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_162_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11002__A1 _00725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09746__A2 _01310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07757__A1 as2650.stack\[11\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09984_ _04001_ _04000_ _04138_ _04140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_89_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_5108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08935_ _03107_ _03177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_130_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11305__A2 _05297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08866_ _03077_ _03112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_111_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07861__I _02250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07817_ _02224_ _02225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_6_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08797_ _03044_ _03041_ _03045_ _03046_ _00208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__11383__I _05455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11069__A1 as2650.stack\[1\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07748_ as2650.stack\[11\]\[2\] _02149_ _02166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11069__B2 as2650.stack\[3\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07679_ _02101_ _02102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09682__A1 _02849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08485__A2 _00615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09788__I _00641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09418_ _03600_ _03601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_90_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10690_ _04397_ _00895_ _04570_ _04798_ _04799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_13_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_185_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08237__A2 _00615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09349_ _02644_ _03548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_142_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06248__A1 _00679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06799__A2 _01239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07996__A1 as2650.stack\[14\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11311_ _05402_ _05403_ _05404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_180_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_180_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12015__CLK clknet_leaf_100_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11242_ _05333_ _05336_ _05265_ _05337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_84_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09737__A2 _01322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07748__A1 as2650.stack\[11\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11544__A2 _00861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11173_ as2650.stack\[14\]\[2\] _05268_ _05269_ as2650.stack\[12\]\[2\] _05215_ _05270_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_121_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06161__B _00619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09028__I _03258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10124_ _03769_ _04272_ _04274_ _04275_ _04276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_164_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_5631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10055_ net40 _04209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_5664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08867__I _03079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07771__I _02128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08173__A1 _02323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_5686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11507__B _03779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07920__A1 _02122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11226__C _03859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09673__A1 _03721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08476__A2 _00886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10957_ _05057_ _05058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_147_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06487__A1 _00928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10283__A2 _01345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10888_ _04752_ _04979_ _04991_ _04992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__10822__A4 _04927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11242__B _05265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11232__A1 _01599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07987__A1 _00728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_1617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11509_ _01992_ _05557_ _05558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_195_1639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_160_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09728__A2 _01254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07739__A1 _02151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08270__C _02578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11535__A2 _02770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08400__A2 _02681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06411__A1 _00833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06981_ _01401_ _01411_ _01418_ _01420_ _01094_ _01421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XTAP_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06962__A2 _01235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05932_ _05757_ _05763_ _05770_ _05785_ _05786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XANTENNA__11299__A1 _02861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08720_ _02456_ _02712_ _02979_ _02987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xclkbuf_leaf_47_wb_clk_i clknet_4_13_0_wb_clk_i clknet_leaf_47_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08777__I _02473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07681__I _02035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_132_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07211__I0 as2650.r123\[0\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08651_ _02918_ _02919_ _02922_ _02923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05863_ as2650.ins_reg\[1\] _05705_ _05717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__09900__A2 _04056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06714__A2 _01155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07602_ _02029_ _02030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_130_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08582_ _02854_ _02855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06297__I _00748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07533_ as2650.stack\[5\]\[14\] _01961_ _01962_ as2650.stack\[4\]\[14\] _01963_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_81_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09664__A1 _02582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06478__A1 _00491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10274__A2 _00822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11471__A1 _00461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07464_ as2650.stack\[9\]\[11\] _01869_ _01758_ as2650.stack\[8\]\[11\] as2650.stack\[10\]\[11\]
+ _01747_ _01897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_62_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09203_ _03418_ _03422_ _03423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06415_ _00860_ _00861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09416__A1 _00677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07395_ _01829_ _01830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_194_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09134_ _03320_ _03323_ _03356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12038__CLK clknet_leaf_15_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_148_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06346_ _00474_ _00586_ _00684_ _00791_ _00512_ _00795_ _00796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai33_1
XANTENNA__09967__A2 _01695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09065_ _01975_ _03252_ _03290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_147_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06277_ _00730_ _00731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_147_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07856__I _01988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09049__S _03271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08016_ _02102_ _02373_ _02377_ _02378_ _00095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__09719__A2 _03875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06760__I _01136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11378__I _05460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10282__I _04418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06402__A1 _00842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09967_ _04075_ _01695_ _04123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08918_ _03069_ _03160_ _03161_ _03162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_150_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09898_ _04049_ _04055_ _04056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_98_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08849_ _03065_ _03096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10231__B _04379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07902__A1 as2650.stack\[10\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11860_ _00229_ clknet_leaf_30_wb_clk_i as2650.r123_2\[0\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10811_ _02194_ _04881_ _04917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_11791_ _00174_ clknet_leaf_84_wb_clk_i as2650.stack\[1\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_2_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09655__A1 _03816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08458__A2 _02722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06469__A1 _00465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10742_ _04847_ _04848_ _04849_ _04797_ _04850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_14_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09311__I _02631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10670__C1 as2650.stack\[10\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10673_ as2650.stack\[13\]\[4\] _01750_ _01755_ as2650.stack\[12\]\[4\] _04783_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__09407__A1 as2650.stack\[6\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09958__A2 _03976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07969__A1 _02334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09467__B _03612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10973__B1 _05057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11225_ _03948_ _01445_ _05202_ _05320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_141_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_1694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10725__B1 _01825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09430__I1 _03285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08394__A1 _02680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11156_ _01150_ _02866_ _03653_ _02851_ _05253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_150_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10107_ _04217_ _04231_ _04260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11087_ _05152_ _05169_ _05184_ _05185_ _05186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_49_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08146__A1 _02323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10038_ _04078_ _04192_ _03727_ _04193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_97_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09894__A1 _04001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_166_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09646__A1 _03794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11989_ _00358_ clknet_leaf_75_wb_clk_i net71 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_182_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11453__A1 _01932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06200_ _00486_ _00505_ _00614_ _00658_ _00659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_31_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11205__A1 as2650.stack\[2\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06880__A1 _01319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07180_ _01565_ _01011_ _01591_ _01299_ _01593_ _01426_ _01618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XANTENNA__09949__A2 _04103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11205__B2 as2650.stack\[0\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_125_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_173_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06131_ _00589_ _00590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_145_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09377__B _03543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06632__A1 _01059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06580__I _00937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06062_ _00520_ _00521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_145_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_195_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11508__A2 _01876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09421__I1 _03261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08385__A1 as2650.stack\[2\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09821_ _03978_ _01428_ _03980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10192__A1 _00601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06935__A2 _01361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09752_ _00731_ _03782_ _03905_ _03912_ _03913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_06964_ _01403_ _01186_ _01230_ _01235_ _01181_ _01404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_100_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08703_ _02705_ _02974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05915_ _05766_ _05726_ _05767_ _05718_ _05768_ _05707_ _05769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_104_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09683_ _03843_ _03844_ _03845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06895_ _01230_ _01235_ _01242_ _01336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_95_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09885__A1 _04041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05846_ _05699_ _05700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08634_ _01732_ _02906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_94_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07360__A2 _01739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08565_ _02834_ _02835_ _05793_ _02837_ _02838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_35_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10247__A2 _04392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07516_ as2650.stack\[9\]\[13\] _01942_ _01941_ as2650.stack\[8\]\[13\] as2650.stack\[11\]\[13\]
+ _01940_ _01947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_08496_ _02730_ _02341_ _02769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_165_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07447_ _01784_ _01878_ _01880_ _01881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_167_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06466__A4 _00615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06871__A1 _01310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07378_ as2650.stack\[7\]\[9\] _01811_ _01812_ as2650.stack\[6\]\[9\] _01813_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_195_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_148_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09117_ _03339_ _03340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06329_ _00778_ _00779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_163_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_178_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09048_ _03162_ _03245_ _03248_ _03275_ _03276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_135_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_163_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07179__A2 _01596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11010_ _02746_ _00502_ _03638_ _05108_ _05109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_145_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10183__A1 net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_161_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output52_I net52 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08128__A1 _01933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05834__I as2650.ins_reg\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_4034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08210__I _02236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_180_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_57_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09876__A1 _01609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11132__B1 _02002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09750__B _03776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11912_ _00281_ clknet_leaf_68_wb_clk_i as2650.ivec\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11843_ _00226_ clknet_leaf_104_wb_clk_i as2650.stack\[7\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_95 io_oeb[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_96_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11435__A1 _00640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06665__I _01108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11774_ _00157_ clknet_leaf_82_wb_clk_i as2650.stack\[3\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08300__A1 _01459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10187__I net91 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_186_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10725_ as2650.stack\[13\]\[5\] _01828_ _01825_ as2650.stack\[12\]\[5\] _04834_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_1997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09976__I net37 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_146_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10656_ _04763_ _04721_ _04764_ _04765_ _04766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_173_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09909__C _03786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11199__B1 _05163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08813__C _03059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10587_ _04533_ _04650_ _04680_ _04698_ _04643_ _04699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_182_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10410__A2 _00704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_108_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_170_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08367__A1 as2650.stack\[3\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11208_ as2650.stack\[1\]\[3\] _05302_ _05303_ as2650.stack\[3\]\[3\] _05304_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__10174__A1 _03684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11139_ _03974_ _05236_ _00360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08119__A1 as2650.stack\[0\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07590__A2 _02015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07327__C1 _01762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_4_2_0_wb_clk_i_I clknet_3_1_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06680_ _00960_ _01121_ _01123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_92_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09619__A1 _03775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10229__A2 _02333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08350_ _02650_ _02651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06575__I _01018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11426__A1 as2650.stack\[9\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_189_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07301_ _01736_ _01737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08281_ _00850_ _02589_ _02590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_162_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_177_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07232_ _01662_ _01668_ _01669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_144_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08790__I _02473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05900__I0 as2650.r123\[2\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11720__CLK clknet_leaf_5_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07163_ _01600_ _01601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06605__A1 _01034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06114_ _00549_ as2650.cycle\[7\] _00573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_121_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10401__A2 _04514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07094_ _01505_ _01528_ _01532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_146_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06045_ _00455_ _00503_ _00504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11870__CLK clknet_leaf_38_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_62_wb_clk_i clknet_4_14_0_wb_clk_i clknet_leaf_62_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_114_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08358__A1 _02516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07030__A1 _01462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09804_ _03933_ _03963_ _03964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_59_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07996_ as2650.stack\[14\]\[1\] _02362_ _02363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_87_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07581__A2 _02006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09735_ _01272_ _01281_ _01283_ _01285_ _03896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_101_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08030__I _02389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06947_ _01372_ _01386_ _01387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_101_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09858__A1 _03925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10468__A2 _03722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09666_ _03818_ _03823_ _03826_ _03827_ _03828_ _03829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_39_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06878_ _01318_ _01319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_83_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08530__A1 _01776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07333__A2 net73 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08617_ _02889_ _02890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_15_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05829_ as2650.ins_reg\[0\] _05683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__11605__B _05647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09597_ _03760_ _03761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_131_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05895__A2 _05748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11417__A1 as2650.stack\[9\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08548_ _01210_ _01135_ _01021_ _02820_ _02821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XANTENNA__11324__C _03813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08479_ _02566_ _02751_ _02752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_71_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10510_ as2650.stack\[7\]\[1\] _01835_ _01790_ as2650.stack\[5\]\[1\] _04623_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_11490_ as2650.r123\[3\]\[2\] _05547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10640__A2 _04704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10441_ _03722_ _04076_ _04555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_164_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05829__I as2650.ins_reg\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08597__A1 _02867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10372_ _03261_ _04490_ _04492_ _04493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_109_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_163_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_105_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08349__A1 _02133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12042_ _00411_ clknet_opt_1_0_wb_clk_i net59 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_3_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10156__A1 _00906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09010__A2 _02495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10470__I _00800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09849__A1 _00800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06609__B _01052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_178_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11408__A1 _03550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05886__A2 _05737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11826_ _00209_ clknet_leaf_106_wb_clk_i as2650.stack\[8\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11743__CLK clknet_leaf_114_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07088__A1 _01520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08285__B1 _02567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11757_ _00140_ clknet_leaf_80_wb_clk_i as2650.stack\[6\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10708_ _00522_ _04800_ _04816_ _04109_ _04817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_105_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11688_ _00071_ clknet_leaf_2_wb_clk_i as2650.stack\[10\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_174_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10639_ _04748_ _04749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__10919__B1 _05007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08115__I _02096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10395__A1 _03609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09001__A2 _03233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11344__B1 _01962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11344__C2 _05180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07850_ _02053_ _02237_ _02248_ _02047_ _00059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_111_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08760__A1 _02461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06801_ _01180_ _01188_ _01238_ _01243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_99_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_85_wb_clk_i_I clknet_4_2_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07781_ net88 _02193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_83_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xinput3 io_in[12] net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_37_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09520_ _00442_ _00782_ _02737_ _03672_ _03684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_49_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06732_ _01168_ _01170_ _01173_ _01174_ _01175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_37_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08785__I _02077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06118__A3 _00576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06663_ _01106_ _01107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_149_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09451_ _02074_ _03617_ _03621_ _03624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_65_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08402_ _02688_ _02689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_91_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06594_ _00489_ _01037_ _01038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10870__A2 net64 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09382_ _03571_ _03562_ _03572_ _03573_ _00266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__09068__A2 _03259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08333_ as2650.stack\[4\]\[11\] _02636_ _02638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_16_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08815__A2 _01131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_177_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08264_ _00686_ _02572_ _02573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_32_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10622__A2 _01839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08291__A3 _02597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07215_ _01546_ _01645_ _01651_ _01652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_08195_ _02213_ _02516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07146_ _01580_ _01583_ _01584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_119_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08025__I _02255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_192_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10386__A1 _03279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07077_ _01515_ _01516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_106_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_156_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_161_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07864__I _02250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06028_ as2650.prefixed _00487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_121_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10138__A1 _02225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07003__A1 _01309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10290__I _04425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09543__A3 _03645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07554__A2 _01910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08751__A1 _02402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06762__B1 _01204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07979_ _02012_ _02348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_19_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08909__B _03079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09718_ _03876_ _02808_ _03879_ _03880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_10990_ _04863_ _05089_ _03737_ _05090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_99_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11335__B _05416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09649_ _03793_ _03809_ _03810_ _03811_ _00552_ _03812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__10310__A1 _01927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07857__A3 _02254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05868__A2 _05721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11611_ _04437_ _05575_ _05647_ _05653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_169_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08806__A2 _00651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08644__B _01733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10893__C _03832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06817__A1 _01257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_54_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11542_ _01773_ _02153_ _05589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_141_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07490__A1 as2650.stack\[14\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11473_ _04525_ _05533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__07490__B2 as2650.stack\[12\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10424_ as2650.stack\[5\]\[0\] _02784_ _02794_ as2650.stack\[4\]\[0\] _04538_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_167_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10377__A1 _03267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06045__A2 _00503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10355_ _00639_ _04375_ _04477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_98_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07774__I _02132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08990__A1 _02368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10129__A1 _02216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10286_ _04422_ _04423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12025_ _00394_ clknet_leaf_39_wb_clk_i as2650.r123\[2\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_111_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11629__A1 net74 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_2_wb_clk_i_I clknet_4_1_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10301__A1 as2650.holding_reg\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_146_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09430__S _03604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11809_ _00192_ clknet_leaf_5_wb_clk_i as2650.stack\[15\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10604__A2 _00896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09470__A2 _00758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07481__B2 as2650.stack\[6\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07000_ _01307_ _01439_ _01440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_174_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11639__CLK clknet_leaf_37_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06036__A2 _00494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_170_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_153_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11580__A3 _01421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08951_ _03115_ _03192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_174_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07902_ as2650.stack\[10\]\[3\] _02274_ _02290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_130_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08882_ _01195_ _03127_ _03128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09525__A3 _01712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07536__A2 _01944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11789__CLK clknet_4_2_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07833_ _02222_ _02237_ _02238_ _02201_ _00052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_56_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07764_ _02177_ _02178_ _02140_ _02179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09503_ _00901_ _02555_ _03667_ _03668_ _03669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
X_06715_ _01120_ _01156_ _01157_ _01158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_112_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11096__A2 _04638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07695_ _01598_ _02084_ _02117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_1642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09434_ _03610_ _00281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06646_ _05695_ _01090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_1664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08500__A4 _02337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09365_ _03558_ _03544_ _03559_ _03560_ _00262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06577_ _01020_ _01021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_21_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07859__I _02256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08316_ _00678_ _02625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_138_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09296_ _03037_ _03494_ _03506_ _03507_ _00246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_55_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09461__A2 _02536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08247_ _00459_ _00798_ _00658_ _02555_ _02556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_20_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08178_ as2650.stack\[7\]\[13\] _02497_ _02503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09213__A2 _03298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07224__A1 as2650.holding_reg\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06027__A2 _00485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07129_ _01565_ _01486_ _01566_ _01567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__11020__A2 _00904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10140_ _04291_ _04280_ _04282_ _04292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_79_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10071_ _00982_ _04225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_43_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07527__A2 _01910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08724__A1 _02989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11991__D _00360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07543__B _01972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05842__I _05688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09314__I _03520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11087__A2 _05169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10973_ _01953_ _04995_ _05057_ _03667_ _05073_ _05074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__06159__B _00617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_44_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10834__A2 _04934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_186_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_175_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_178_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_157_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09452__A2 _03613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_156_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07463__A1 _01894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11525_ _02625_ _05573_ _05574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_106_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_172_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11456_ _01622_ _05498_ _05513_ as2650.r123\[2\]\[6\] _05518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_156_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09204__A2 _03423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10407_ _00519_ _00893_ _00565_ _04311_ _04521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_125_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11011__A2 _02759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11387_ _02678_ _05457_ _05461_ _05466_ _00378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__06622__B _01021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06569__A3 _00983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07766__A2 _02163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_180_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11931__CLK clknet_leaf_62_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10338_ _04464_ _00331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_113_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10770__A1 _04875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_119_wb_clk_i clknet_4_2_0_wb_clk_i clknet_leaf_119_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_191_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10269_ _03712_ _04320_ _04407_ _04408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_113_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07518__A2 _01812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08715__A1 as2650.stack\[15\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12008_ _00377_ clknet_leaf_117_wb_clk_i as2650.stack\[9\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_78_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10522__A1 as2650.stack\[13\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08549__B _02590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10522__B2 as2650.stack\[12\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10798__C _04904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06848__I _01103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09140__A1 _05759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06500_ _00943_ _00944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07480_ _01836_ _01912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_34_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10825__A2 _04930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09691__A2 _03849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06431_ _00617_ _00869_ _00875_ _00876_ _00877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_179_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07679__I _02101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09150_ _03314_ _03348_ _03371_ _03372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_148_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09979__B1 _04134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06362_ _00808_ _00809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_159_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09443__A2 _03617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_187_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08101_ _02439_ _02445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09081_ _01569_ _01204_ _01637_ _03304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_06293_ _00744_ _00745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_120_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11250__A2 _05344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08032_ _02250_ _02392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_162_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_190_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07206__A1 as2650.r0\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11002__A2 _00866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07757__A2 _02149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08954__A1 _01602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09983_ _02125_ _04136_ _04051_ _04138_ _04139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_89_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10761__A1 _04237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08934_ as2650.r123_2\[1\]\[5\] _03105_ _03176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_131_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_192_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09843__B _04001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10989__B _04332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08865_ _03057_ _03111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_29_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07816_ net68 _02224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_79_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06193__A1 _00460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08796_ as2650.stack\[8\]\[5\] _03035_ _03021_ _03046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_85_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07747_ _02051_ _02141_ _02162_ _02165_ _00039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__11069__A2 _05162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07678_ _02100_ _02101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09682__A2 _01261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09417_ _03598_ _03599_ _03600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06629_ _01068_ _01070_ _01072_ _01073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_129_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11613__B _04441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11804__CLK clknet_leaf_3_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06493__I _00936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09348_ as2650.stack\[3\]\[0\] _03546_ _03547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_179_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06248__A2 _00574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09279_ _03493_ _03494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_166_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07996__A2 _02362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11310_ as2650.stack\[10\]\[6\] _05180_ _05269_ as2650.stack\[8\]\[6\] _05174_ _05403_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_148_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11241_ _05334_ _05335_ _05336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_88_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07748__A2 _02149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11544__A3 _05589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11172_ _01900_ _05269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10752__A1 _04811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10123_ _03991_ _04275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_122_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10054_ _04129_ _04204_ _04207_ _04024_ _04208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_121_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10504__A1 _04610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08173__A2 _02489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09370__A1 _03561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06668__I _01111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06184__A1 _00639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07920__A2 _02292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05931__A1 _05771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_4_7_0_wb_clk_i_I clknet_3_3_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10956_ _05056_ _05057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08476__A3 _02598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06487__A2 _00930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11523__B _05539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10887_ _03816_ _04978_ _04363_ _04991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_31_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11232__A2 _05140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09928__B _03761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_160_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11508_ _01990_ _01876_ _05557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05998__A1 _05720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10991__A1 _03816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11439_ _05496_ _03374_ _05506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07448__B _01881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09728__A3 _01258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_47_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_153_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_154_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06980_ _01390_ _00764_ _01419_ _01420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07962__I _05671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input6_I io_in[34] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05931_ _05771_ _05773_ _05779_ _05784_ _05785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_117_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09361__A1 _03555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07211__I1 as2650.r123_2\[0\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06578__I _01021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08650_ _01764_ _02920_ _02921_ _02922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_05862_ _05708_ _05715_ _05716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06175__A1 as2650.cycle\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07601_ _02027_ _02028_ _02029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_94_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08581_ _02853_ _02854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_81_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11827__CLK clknet_leaf_106_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07532_ _01827_ _01962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_81_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_165_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_16_wb_clk_i clknet_4_4_0_wb_clk_i clknet_leaf_16_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_1_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09664__A2 _00815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06478__A2 _00898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10828__I _04922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07463_ _01894_ _01895_ _01846_ _01896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__07675__A1 as2650.stack\[13\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11471__A2 _00493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09202_ _03420_ _03421_ _03422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_06414_ _00843_ _00859_ _00860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_10_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_195_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07394_ _01828_ _01829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09416__A2 _00921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09133_ _03353_ _03325_ _03354_ _03355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07427__A1 _01854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06345_ _00794_ _00795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__11223__A2 _05318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09064_ _03284_ _03288_ _03289_ _00232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_120_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06276_ _00729_ _00730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10982__A1 _02235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08015_ as2650.stack\[14\]\[5\] _02360_ _02356_ _02378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_163_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08927__A1 _01430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10734__A1 _02107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06402__A2 _00847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09966_ _04116_ _04121_ _04122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_104_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08917_ _01350_ _03096_ _03161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_103_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09897_ _04013_ _03999_ _04051_ _04055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_24_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08848_ _03071_ _03091_ _03094_ _03095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_4249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07902__A2 _02274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08779_ _03028_ _03022_ _03030_ _03032_ _00204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_2825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09104__A1 as2650.r0\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09799__I _03879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10810_ _04595_ _04916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11790_ _00173_ clknet_leaf_84_wb_clk_i as2650.stack\[1\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08458__A3 _01037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10741_ _01465_ _05737_ _04849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10738__I _04844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_144_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10670__B1 _01817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_35_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10670__C2 _01875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10672_ as2650.stack\[15\]\[4\] _02781_ _01779_ as2650.stack\[14\]\[4\] _04782_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__11062__C _05160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09407__A2 _03585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_142_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07969__A2 _02337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10973__A1 _01953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10973__B2 _03667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10473__I _00698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11224_ _04275_ _01429_ _05319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_135_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10725__A1 as2650.stack\[13\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10725__B2 as2650.stack\[12\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08394__A2 _02681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11155_ _01269_ _05241_ _05248_ _05251_ _05252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_96_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10106_ _02218_ _04101_ _04258_ _04259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_5440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11086_ _00755_ _05185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_5451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08146__A2 _02468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10037_ _04169_ _04191_ _04192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_64_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11237__C _05174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11150__A1 net49 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09894__A2 _04000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11988_ _00357_ clknet_leaf_70_wb_clk_i net69 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_90_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10939_ _02224_ _05040_ _05041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_177_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06347__B _00796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_140_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11205__A2 _05296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06130_ _05771_ _00589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10964__A1 _02229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_134_wb_clk_i clknet_4_1_0_wb_clk_i clknet_leaf_134_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_69_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06061_ _00519_ _00520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_195_1459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_160_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_132_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08909__A1 _03150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10716__A1 _02906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09820_ _03978_ _01428_ _03979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_140_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10192__A2 _04341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09751_ _03908_ _03910_ _03911_ _03912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06963_ _01179_ _01403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_100_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08702_ as2650.stack\[15\]\[0\] _02972_ _02973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09334__A1 as2650.stack\[4\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05914_ as2650.r123\[1\]\[3\] as2650.r123\[0\]\[3\] as2650.r123_2\[1\]\[3\] as2650.r123_2\[0\]\[3\]
+ _05683_ _05712_ _05768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_80_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09682_ _02849_ _01261_ _03844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06148__A1 _00601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06894_ _01334_ _01335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_82_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08633_ _02897_ _02904_ _00647_ _02905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05845_ as2650.ins_reg\[4\] _05699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_110_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08564_ _02836_ _02837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_74_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_120_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07515_ _01943_ _01945_ _01799_ _01946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08495_ _02583_ _02768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_145_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07446_ as2650.stack\[13\]\[10\] _01816_ _01879_ as2650.stack\[12\]\[10\] _01880_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08028__I _02387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06320__A1 _00763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07377_ _01781_ _01812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_136_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09116_ _00640_ _03103_ _03338_ _03339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_149_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06328_ _00513_ _00778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08073__A1 _02314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10955__A1 net69 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11389__I _05460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09047_ _03273_ _03262_ _03274_ _03275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07820__A1 as2650.stack\[14\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06259_ _00714_ _00632_ _00715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_135_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10707__A1 _00521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_150_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08698__I _02709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06387__A1 _00825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10183__A2 _04333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09949_ _03866_ _04103_ _04104_ _04087_ _04105_ _04106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_150_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09325__A1 _02449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11132__A1 as2650.stack\[14\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output45_I net45 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09876__A2 _01596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06011__I _00469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11911_ _00280_ clknet_leaf_71_wb_clk_i as2650.ivec\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_4079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_185_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08647__B _01764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11842_ _00225_ clknet_leaf_102_wb_clk_i as2650.stack\[7\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_36_wb_clk_i_I clknet_4_6_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09628__A2 _03790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05850__I _05700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_96 io_oeb[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_1943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11435__A2 _01106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11773_ _00156_ clknet_leaf_91_wb_clk_i as2650.stack\[4\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07103__A3 _01517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08300__A2 _02608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10724_ as2650.stack\[15\]\[5\] _04822_ _01822_ as2650.stack\[14\]\[5\] _04833_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_159_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10655_ _01434_ _05761_ _04765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__11199__A1 as2650.stack\[5\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08382__B _02671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11199__B2 as2650.stack\[7\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08064__A1 _02302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10586_ _04620_ _04649_ _04697_ _04640_ _04698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_155_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10946__A1 _04226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10136__C _01291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_190_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11672__CLK clknet_leaf_131_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11207_ _01863_ _05303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08367__A2 _02645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11138_ _03261_ _05189_ _05208_ _05235_ _05236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_96_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_75_wb_clk_i_I clknet_4_11_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08119__A2 _02445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11069_ as2650.stack\[1\]\[0\] _05162_ _05163_ as2650.stack\[3\]\[0\] _05167_ _05168_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XTAP_5281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07327__B1 _01761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09433__S _03600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_188_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06856__I _00437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06550__A1 _00532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_51_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11426__A2 _05476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07300_ _01730_ _01736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_149_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08280_ _00873_ _02589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_149_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06302__A1 _00662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07231_ _01666_ _01667_ _01668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06853__A2 _01249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10237__I0 _02845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07687__I _02109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07162_ _05716_ _05722_ _05729_ _01600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__08055__A1 as2650.stack\[12\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10937__A1 _04590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10327__B _00507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06113_ _00485_ _00571_ _00572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07093_ _00999_ _01502_ _01531_ _00019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_12_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06044_ _05699_ _00503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_105_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09803_ _03906_ _03962_ _03963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_114_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07995_ _02359_ _02362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_87_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09307__A1 _03047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09734_ _01281_ _01283_ _01285_ _01273_ _03895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_99_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06946_ _01367_ _01385_ _01386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_28_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_31_wb_clk_i clknet_4_7_0_wb_clk_i clknet_leaf_31_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_132_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09858__A2 _04011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09665_ _02332_ _03752_ _03787_ _03828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06877_ _01016_ _00977_ _01318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_27_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08616_ _01711_ _02889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_27_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05828_ net94 _05682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_82_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09596_ _00722_ _03760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_131_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_128_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08547_ _01597_ _01459_ _01430_ _01265_ _02820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XANTENNA__10288__I _04424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11417__A2 _05476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08981__I _03219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08294__A1 _02594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08478_ _02577_ _02750_ _02751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07429_ _01795_ _01863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_137_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06715__B _01157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07597__I _02024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08046__A1 as2650.stack\[12\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10440_ _03665_ _04554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_109_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10928__A1 _05026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09794__A1 _03951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11695__CLK clknet_leaf_120_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10371_ _03138_ _04491_ _04492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_139_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09518__S _03682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_156_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11994__D _00363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_191_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08349__A2 _02649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09546__A1 _03707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12041_ _00410_ clknet_leaf_9_wb_clk_i net70 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_137_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_172_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10156__A2 _00986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05845__I as2650.ins_reg\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11353__A1 _02347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08221__I _02529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07265__C _00943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11105__A1 _03948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06780__A1 _01202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09849__A2 _02618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_189_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06676__I _01118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10864__B1 _04947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09052__I _01927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10198__I _03875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11825_ _00208_ clknet_leaf_100_wb_clk_i as2650.stack\[8\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11408__A2 _05473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07088__A2 _01526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08285__A1 _02592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11756_ _00139_ clknet_leaf_80_wb_clk_i as2650.stack\[6\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_186_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08285__B2 _01038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10092__A1 _04129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10707_ _00521_ _04807_ _04813_ _04815_ _04816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__10092__B2 _04024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11687_ _00070_ clknet_leaf_126_wb_clk_i as2650.stack\[10\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_144_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10638_ _04747_ _04748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_155_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10147__B _04298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10919__A1 _01904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10919__B2 _03667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10569_ _01744_ _04681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_143_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11592__A1 net49 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09428__S _03604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_170_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09537__A1 _02594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10661__I _04332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11344__A1 as2650.stack\[8\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11344__B2 as2650.stack\[11\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07175__C _01027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06800_ _01180_ _01188_ _01237_ _01242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_96_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08760__A2 _02695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07780_ _02084_ _02192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_42_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput4 io_in[13] net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_110_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06731_ _01169_ _00665_ _01174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_37_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09450_ as2650.stack\[5\]\[2\] _03615_ _03623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06662_ _01105_ _01106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_64_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06586__I net78 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06523__A1 _00963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08401_ _02030_ _02649_ _02664_ _02688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_1857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_149_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09381_ _02129_ _02653_ _03543_ _03573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06593_ _00596_ _01037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_51_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08332_ _02516_ _02628_ _02633_ _02637_ _00152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_33_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06826__A2 _01267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08263_ _00645_ _00747_ _02572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_18_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07214_ _01646_ _01647_ _01650_ _01651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_119_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08194_ _02513_ _02508_ _02512_ _02515_ _00136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_158_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09776__A1 _03933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07145_ _01491_ _01410_ _01581_ _01582_ _01583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_180_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_145_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07076_ as2650.r123\[0\]\[5\] as2650.r123_2\[0\]\[5\] _05710_ _01515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07251__A2 _01687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06027_ _00483_ _00485_ _00486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_161_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10138__A2 _04101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11335__A1 _05796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07003__A2 _01284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08200__A1 as2650.stack\[6\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08041__I _02066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08751__A2 _02996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07978_ _02346_ _02347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06762__A1 _01203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07880__I _01762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06762__B2 _01101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09717_ _03752_ _03878_ _03879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06929_ _01352_ _01369_ _01370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__11616__B _05647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07813__C _02210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09648_ _03771_ _03811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06496__I _05714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06514__A1 _00663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10310__A2 _04439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09579_ _00681_ _03743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_167_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11610_ _00697_ _05652_ _00415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_73_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08267__A1 _05698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11541_ _04460_ _05575_ _05571_ _05540_ _05588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__06817__A2 _01123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_128_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08019__A1 _02113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11472_ _05530_ _05531_ _05532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07490__A2 _01877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_167_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09767__A1 _02082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10423_ as2650.stack\[7\]\[0\] _04536_ _01744_ as2650.stack\[6\]\[0\] _04537_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__09767__B2 _03878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11574__A1 _00427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10354_ _00715_ _00906_ _04310_ _04475_ _04476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_152_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09519__A1 _02625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08990__A2 _02500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10285_ _04419_ _04421_ _00966_ _00911_ _04422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_97_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10129__A2 _01609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11326__A1 net77 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12024_ _00393_ clknet_leaf_35_wb_clk_i as2650.r123\[2\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_78_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09534__A4 _03697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07790__I _02187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06505__A1 _00948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10301__A2 _04423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_185_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_178_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08258__A1 _00557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11808_ _00191_ clknet_leaf_5_wb_clk_i as2650.stack\[15\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_61_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_147_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06808__A2 _00987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11739_ _00122_ clknet_leaf_113_wb_clk_i as2650.stack\[8\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06355__B _00803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07481__A2 _01912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07965__I _02333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11565__A1 _02965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08950_ as2650.r123_2\[1\]\[6\] _03105_ _03191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_131_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11317__A1 _05185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07901_ _02067_ _02270_ _02288_ _02289_ _00069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_69_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08881_ _03065_ _03127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_130_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09525__A4 _02580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07832_ as2650.stack\[14\]\[14\] _02188_ _02238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_61_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_135_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07763_ _02155_ _02178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_96_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09502_ _00825_ _02352_ _00648_ _03668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06714_ _00976_ _01155_ _01157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_96_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08497__A1 _02348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07694_ _02115_ _02116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_129_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09433_ as2650.ivec\[6\] _03609_ _03600_ _03610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06645_ _01086_ _01069_ _01084_ _01088_ _01089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_53_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_59_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_169_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09364_ _03231_ _03548_ _03553_ _03560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_52_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_75_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06576_ _05776_ _01020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_24_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_80_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10056__A1 net39 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08315_ _02610_ _02605_ _02624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_127_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09997__A1 _03734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09295_ _03231_ _02673_ _03500_ _03507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_36_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09049__I0 _03276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08246_ _02554_ _02555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_36_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08177_ _02325_ _02500_ _02501_ _02502_ _00132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_192_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11556__A1 _00736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07128_ as2650.holding_reg\[6\] _00829_ _01566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_137_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07224__A2 _01486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08421__A1 as2650.stack\[1\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07775__A3 _02034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07059_ _01088_ _01498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_106_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06983__A1 _00430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11733__CLK clknet_leaf_111_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10070_ _04199_ _03871_ _04211_ _00688_ _00817_ net40 _04224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai222_2
XFILLER_134_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_102_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08724__A2 _02712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10531__A2 _04582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10972_ _00522_ _05059_ _05072_ _05073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_56_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08488__A1 _02758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10295__A1 as2650.holding_reg\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_169_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09330__I _02632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10047__A1 _04175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09988__A1 _00633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11244__B1 _05269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11524_ _05569_ _02001_ _05572_ _05573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_102_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11455_ _02089_ _00866_ _00657_ _03100_ _05517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_137_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11547__A1 _02027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07785__I _02196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10406_ _04411_ _04520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_124_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11386_ as2650.stack\[9\]\[11\] _05464_ _05466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_139_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08963__A2 _03203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10337_ _04462_ _04463_ _04457_ _00781_ _04464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_139_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06974__A1 _01392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_136_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10268_ _02569_ _02964_ _04406_ _04407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_140_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12007_ _00376_ clknet_4_2_0_wb_clk_i as2650.stack\[9\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08715__A2 _02972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10199_ _02572_ _04349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10522__A2 _01829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11256__B _00914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08479__A1 _02566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07025__I net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07151__A1 _01166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_179_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06430_ _00543_ _00867_ _00876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_2090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_146_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10038__A1 _04078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09979__A1 _00719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09979__B2 _03995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06361_ _00627_ _00808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_33_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08100_ _02060_ _02430_ _02444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_124_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09080_ _03301_ _03302_ _03303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_175_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06292_ _00743_ _00528_ _00744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_147_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08031_ as2650.stack\[12\]\[0\] _02390_ _02391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11538__A1 _05556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11538__B2 _04298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07206__A2 _01216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11756__CLK clknet_leaf_80_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11002__A3 _03766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10210__A1 net91 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09982_ _04046_ _04048_ _04092_ _04138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_88_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout94_I net53 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06965__A1 _01342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10761__A2 _04866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08933_ _03110_ _03174_ _03175_ _00215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_118_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08864_ _03068_ _03110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_170_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05943__I _05749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07815_ _01380_ _02223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_3708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11166__B _05222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05925__C1 _05778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08795_ _02376_ _03029_ _03045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06193__A2 _00454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07746_ as2650.stack\[11\]\[1\] _02163_ _02164_ _02165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_2_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10277__A1 _01008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07677_ net52 _02100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_52_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09416_ _00677_ _00921_ _00883_ _00768_ _03599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_06628_ _01015_ _00828_ _01071_ _01072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11613__C _05185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08890__A1 _00426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10029__A1 _03759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10029__B2 _03811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09347_ _03545_ _03546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_178_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06559_ _00714_ _00555_ _00973_ _01002_ _01003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_166_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06248__A3 _00704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09278_ _02669_ _03493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_154_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06653__B1 _01072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08229_ _02530_ _02541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11529__A1 _02648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_193_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11240_ as2650.stack\[6\]\[4\] _02387_ _02271_ as2650.stack\[4\]\[4\] _05298_ _05335_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_107_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_107_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11171_ _01811_ _05268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_122_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06956__A1 as2650.holding_reg\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10752__A2 _04844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output75_I net75 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10122_ _04270_ _04273_ _04274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_122_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_164_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_164_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07554__B _01982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10053_ _04200_ _04205_ _04206_ _04207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_103_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06708__A1 _01150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10504__A2 _04615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09370__A2 _03562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06184__A2 _00640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_95_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_169_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05931__A2 _05773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10268__A1 _02569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10955_ net69 _05031_ _05056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__07133__A1 _01569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_186_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10886_ _04725_ _04979_ _04988_ _04989_ _04990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_31_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11507_ _00823_ _04554_ _03779_ _05556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_89_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_1608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_156_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05998__A2 _00454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09189__A2 _03405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10991__A2 _05080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11438_ _05497_ _05505_ _00390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09433__I0 as2650.ivec\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09728__A4 _01260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11369_ _05453_ _00373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_28_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09663__C _03825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05930_ _05781_ _05725_ _05782_ _05717_ _05783_ _05706_ _05784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XTAP_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10602__C _04419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05861_ as2650.r123\[1\]\[7\] as2650.r123\[0\]\[7\] as2650.r123_2\[1\]\[7\] as2650.r123_2\[0\]\[7\]
+ _05685_ _05714_ _05715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_120_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_27_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06175__A2 _00632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07600_ _01729_ _02028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_82_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_94_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08580_ _02852_ _02853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_130_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07531_ _01900_ _01961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__11456__B1 _05513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07462_ as2650.stack\[2\]\[11\] _01865_ _01866_ _01895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_62_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08872__A1 _01150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07675__A2 _02062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09201_ _05743_ _01517_ _03421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_165_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06413_ _00831_ _00844_ _00859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__11208__B1 _05303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07393_ _01750_ _01828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_56_wb_clk_i clknet_4_15_0_wb_clk_i clknet_leaf_56_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_124_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09416__A3 _00883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09132_ _03326_ _03330_ _03354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_06344_ _00793_ _00794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_31_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08624__A1 _02347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09063_ as2650.r123_2\[0\]\[5\] _03284_ _03289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_120_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_175_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06275_ _00470_ _00729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_135_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05938__I _05784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08014_ _02376_ _02365_ _02377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09424__I0 as2650.ivec\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_191_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08927__A2 _03111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10734__A2 _04789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09965_ _04118_ _04120_ _04121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_103_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08916_ _03071_ _03158_ _03159_ _03160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_135_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09896_ _03774_ _04053_ _03813_ _04054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_115_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10498__A1 net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08847_ _03092_ _03093_ _03094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08778_ as2650.stack\[8\]\[1\] _03026_ _03031_ _03032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_2804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_26_wb_clk_i_I clknet_4_5_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07729_ _02148_ _02149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07821__C _02210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07115__A1 _05742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_3_3_0_wb_clk_i clknet_0_wb_clk_i clknet_3_3_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__08458__A4 _00834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10740_ _04229_ _05746_ _04848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_25_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10670__A1 as2650.stack\[9\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10670__B2 as2650.stack\[8\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10671_ as2650.stack\[11\]\[4\] _01738_ _01786_ _04781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_179_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08615__A1 _00958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07549__B _01978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_154_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08224__I _02529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11223_ _05281_ _05318_ _00362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_194_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09040__A1 _03267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_162_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10725__A2 _01828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_194_1696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11154_ _03138_ _02815_ _05249_ _05250_ _05241_ _05251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_46_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10105_ _04254_ _04257_ _04258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_133_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_95_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11085_ _05170_ _05183_ _05184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_5441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10036_ _04170_ _04150_ _04191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10489__A1 _04585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11987_ _00356_ clknet_leaf_77_wb_clk_i net68 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_17_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08854__A1 _01103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10938_ _02216_ _02211_ _04949_ _05040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__07303__I _01738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10869_ _04167_ _04789_ _04971_ _04973_ _04912_ _00353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_34_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08606__B2 _01416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_160_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10964__A2 _05064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06060_ _00518_ _00519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08134__I _02470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_173_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07973__I _02341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_103_wb_clk_i clknet_4_9_0_wb_clk_i clknet_leaf_103_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_141_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_86_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06962_ _01230_ _01235_ _01402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09750_ _03908_ _03910_ _03776_ _03911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_101_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_189_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05913_ as2650.r123\[2\]\[3\] as2650.r123_2\[2\]\[3\] _05712_ _05767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_95_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08701_ _02971_ _02972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_171_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09681_ _01254_ _01258_ _01260_ _01273_ _03843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
X_06893_ _01331_ _01333_ _01334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__06148__A2 _00517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08632_ _00958_ _01686_ _02900_ _02903_ _02904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_05844_ _05697_ _05690_ _05698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_54_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08563_ _01565_ _02836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_70_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07514_ as2650.stack\[2\]\[13\] _01944_ _01866_ _01945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08845__A1 _01120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08494_ _02752_ _02763_ _02766_ _02767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__08309__I _02331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_184_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07445_ _01818_ _01879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10652__A1 _02619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06320__A2 _00765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07376_ _01810_ _01811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09115_ _05697_ _03256_ _03338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__10404__A1 _03714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06327_ _00564_ _00690_ _00777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_109_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08073__A2 _02420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06084__A1 _00469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10955__A2 _05031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09046_ _01904_ _03250_ _03274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06258_ _00548_ _00713_ _00714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_136_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07820__A2 _02208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09022__A1 _01800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06189_ _00494_ _00648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_85_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10707__A2 _04807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06720__C _01055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06387__A2 _00832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10183__A3 _03968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09948_ _00957_ _04105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_131_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09325__A2 _03523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09879_ _03987_ _04035_ _04036_ _04037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_57_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11132__A2 _05225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11910_ _00279_ clknet_leaf_70_wb_clk_i as2650.ivec\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_85_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10340__B1 _04343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_161_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output38_I net38 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11841_ _00224_ clknet_leaf_102_wb_clk_i as2650.stack\[7\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_97 io_oeb[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_163_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08836__A1 _01043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08219__I _02534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11772_ _00155_ clknet_leaf_91_wb_clk_i as2650.stack\[4\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_54_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11435__A3 _05502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10643__A1 _04654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10723_ _02789_ _04830_ _04831_ _04832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_109_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10654_ _01434_ _05761_ _04764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_139_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11199__A2 _05162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07279__B _01305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08064__A2 _02258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10585_ _04622_ _04696_ _04697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_139_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10946__A2 _05028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_1_wb_clk_i clknet_4_1_0_wb_clk_i clknet_leaf_1_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_86_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09013__A1 _03243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08889__I _03059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07793__I net87 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11206_ _01870_ _05302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_79_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10174__A3 _04305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11137_ _05220_ _05234_ _05148_ _05235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_190_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11068_ _05166_ _05167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_95_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07327__A1 as2650.stack\[3\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07327__B2 as2650.stack\[0\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08524__B1 _01745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_168_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10019_ _04173_ _04174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_64_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_91_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_52_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06550__A2 _00991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06302__A2 _00608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07968__I _02336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07230_ as2650.holding_reg\[7\] _00871_ _01667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_81_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06805__C _01165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10237__I1 _04157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07161_ _01451_ _01599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_121_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06066__A1 _00523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10937__A2 _05030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06112_ _00570_ _00571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_145_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07092_ as2650.r123\[1\]\[5\] _01197_ _01530_ _01107_ _01531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_145_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06043_ _00501_ _00502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_145_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09004__A1 _03044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11347__C1 as2650.stack\[14\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07566__A1 _01991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09802_ _03838_ _03864_ _03907_ _03918_ _03962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_99_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07994_ _01984_ _02357_ _02358_ _02361_ _00090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_87_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10570__B1 _04681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_190_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_101_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09307__A2 _03508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06945_ _01383_ _01384_ _01385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09733_ _03762_ _03894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07318__A1 net86 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09712__C1 _00818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10997__C _05076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06876_ _01316_ _01298_ _01317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09664_ _02582_ _00815_ _03827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09423__I _03600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08615_ _00958_ _01686_ _02887_ _02888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_05827_ _05680_ _05681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09595_ _00538_ _03759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10569__I _01744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_71_wb_clk_i clknet_4_11_0_wb_clk_i clknet_leaf_71_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_36_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08546_ _02818_ _02819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_42_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_145_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10625__A1 as2650.stack\[11\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08477_ _00898_ _00598_ _00616_ _01130_ _02750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_126_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09491__A1 _03657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07428_ _01739_ _01862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_156_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06844__A3 _01285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07359_ _01794_ _01795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_195_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09243__A1 _03439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_148_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08046__A2 _02390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06057__A1 _00514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10928__A2 _04228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10370_ _04482_ _04491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09029_ _03255_ as2650.r123_2\[0\]\[0\] _03259_ _03260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_108_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12040_ _00409_ clknet_leaf_9_wb_clk_i net73 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_116_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08349__A3 _02254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11105__A2 _01161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06780__A2 _01221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10864__B2 _04534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08809__A1 _01050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11824_ _00207_ clknet_leaf_100_wb_clk_i as2650.stack\[8\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10616__A1 _04609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08285__A2 _02593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09489__B _02761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11755_ _00138_ clknet_leaf_81_wb_clk_i as2650.stack\[6\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06906__B _01346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07788__I _02199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10706_ _04397_ _04723_ _04814_ _04815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_105_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11686_ _00069_ clknet_leaf_124_wb_clk_i as2650.stack\[10\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_146_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10637_ _03958_ _04746_ _04747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_122_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06048__A1 _05675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10568_ _00517_ _04665_ _04679_ _04583_ _04680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_142_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08993__B1 _03227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11592__A2 _05635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_127_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_48_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10499_ _03795_ _05782_ _04612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_114_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09537__A2 _02602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08412__I _02688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11259__B _00847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07548__A1 _01622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08745__B1 _03003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11344__A2 _05226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_68_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput5 io_in[33] net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06730_ _01171_ _01064_ _01172_ _01067_ _01173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XTAP_5090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06661_ _01103_ _00835_ _01104_ _01105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_1814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06523__A2 _00966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08400_ _02686_ _02681_ _02682_ _02687_ _00170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_80_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_149_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09380_ as2650.stack\[3\]\[7\] _03552_ _03572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06592_ _01035_ _01036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10607__A1 _02619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08331_ as2650.stack\[4\]\[10\] _02636_ _02637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_166_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09473__A1 _00622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08276__A2 _01723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06816__B _01257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06287__A1 _00518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11280__A1 as2650.stack\[11\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08262_ _02570_ _02571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_60_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07213_ _05774_ _01649_ _01650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09225__A1 _03439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08193_ as2650.stack\[6\]\[9\] _02514_ _02515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_118_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07144_ _01480_ _01488_ _01582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09776__A2 _03935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_145_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07787__A1 _02198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_161_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07075_ _01511_ _01512_ _01513_ _01514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__10852__I _04946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_192_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09418__I _03600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06026_ _00484_ _00485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05893__S0 _05684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_3_1_0_wb_clk_i_I clknet_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09862__B _03883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06211__A1 _00500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07977_ _02345_ _02346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06762__A2 _01112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10801__B _04907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09716_ _03665_ _03877_ _03878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__11099__A1 _02813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06928_ _01367_ _01368_ _01369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09700__A2 _03790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10846__A1 _04949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09647_ net31 _03773_ _03810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_16_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06859_ _00437_ _01252_ _01300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_16_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06514__A2 _00461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09578_ _03741_ _03742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_82_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08529_ _01787_ _02800_ _02801_ _02802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_93_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09464__A1 _02119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08267__A2 _02570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11271__A1 as2650.stack\[4\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11540_ _02648_ _05576_ _05587_ _00410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_141_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_184_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07401__I _01835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11471_ _00461_ _00493_ _00518_ _02010_ _05531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__08019__A2 _02373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_109_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11023__A1 _05120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12018__CLK clknet_leaf_101_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10422_ _01737_ _04536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09767__A2 _03879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06017__I _05688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_178_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_193_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08975__B1 _03214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11574__A2 _02813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10353_ _03991_ _04307_ _04474_ _04475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_136_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05884__S0 _05684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10284_ _00767_ _04420_ _00765_ _03749_ _04421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_2_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12023_ _00392_ clknet_leaf_38_wb_clk_i as2650.r123\[2\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_133_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06202__A1 _00647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10837__A1 _04937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06505__A2 _00449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07702__A1 as2650.stack\[13\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_178_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11807_ _00190_ clknet_leaf_134_wb_clk_i as2650.stack\[15\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08258__A2 _02004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09455__A1 _03558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06269__A1 _00711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11262__A1 _03149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07466__B1 _01877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11738_ _00121_ clknet_leaf_114_wb_clk_i as2650.stack\[8\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08407__I _02693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06808__A3 _00995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07311__I _01746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11669_ _00052_ clknet_leaf_128_wb_clk_i as2650.stack\[14\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_89_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11014__A1 _03650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11014__B2 _00555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07769__A1 _02113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11565__A2 _05521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06441__A1 _00886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08142__I _02466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_139_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07900_ _02167_ _02285_ _02286_ _02289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_155_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08880_ _03124_ _01127_ _03125_ _03126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_44_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07981__I _02349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08194__A1 _02513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07831_ _02236_ _02237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06597__I net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07762_ _02109_ _02177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05952__B1 _05762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10340__C _04456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09501_ _03666_ _03667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06713_ _00976_ _01155_ _01156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_07693_ net62 _02115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09694__A1 _03819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_168_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_183_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09432_ _01975_ _03609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06644_ _01087_ _01088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_06575_ _01018_ _01019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_146_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09363_ as2650.stack\[3\]\[3\] _03546_ _03559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_181_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10056__A2 net38 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08314_ _02606_ _02622_ _02623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__11253__A1 _03279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09997__A2 _04152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09294_ as2650.stack\[2\]\[3\] _03496_ _03506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_177_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08245_ _00743_ _00925_ _02554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_123_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08176_ as2650.stack\[7\]\[12\] _02497_ _02502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_118_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11556__A2 _02841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07127_ _05797_ _01565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_119_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08421__A2 _02697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07058_ _01485_ _01488_ _01497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_161_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06983__A2 _05808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06009_ as2650.cycle\[0\] _00468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08987__I _02493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10819__A1 _03740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09685__A1 _03842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10971_ _00783_ _05069_ _05071_ _04364_ _04554_ _05072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__08488__A2 _02760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output20_I net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11244__A1 as2650.stack\[14\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11244__B2 as2650.stack\[12\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07131__I _05743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11523_ _04437_ _05570_ _05571_ _05539_ _05572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_11_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_172_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06671__A1 _00695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11454_ _05515_ _05516_ _00395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_7_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_125_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10706__B _04814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08948__B1 _03189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11547__A2 _05579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10405_ _04351_ _04517_ _04518_ _04519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_11385_ _02675_ _05457_ _05461_ _05465_ _00377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_152_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09058__I _03271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06423__A1 _00765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10336_ _00750_ _04463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_152_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10267_ _03673_ _02741_ _03692_ _04406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_171_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12006_ _00375_ clknet_leaf_117_wb_clk_i as2650.stack\[9\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_113_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10198_ _03875_ _04348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_113_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07306__I net48 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09676__A1 net89 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11483__A1 _05264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_opt_1_0_wb_clk_i_I clknet_4_1_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_128_wb_clk_i clknet_4_0_0_wb_clk_i clknet_leaf_128_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_61_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_163_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06360_ _00543_ _00806_ _00807_ _00005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11235__A1 _05813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10038__A2 _04192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09979__A2 _04130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08137__I _02473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08100__A1 _02060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_148_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06291_ as2650.cycle\[6\] _00743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07976__I _01663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08030_ _02389_ _02390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_159_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10616__B _04726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09600__A1 _03740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_4_5_0_wb_clk_i clknet_3_2_0_wb_clk_i clknet_4_5_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_85_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06414__A1 _00843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10210__A2 _00971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09981_ net88 _04136_ _04137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_118_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06965__A2 _01326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08932_ _01387_ _03163_ _03130_ as2650.r123_2\[1\]\[4\] _03175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_170_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout87_I net65 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_130_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08863_ _03068_ _03098_ _03106_ _03109_ _00211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_112_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_85_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06717__A2 _01158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07914__A1 as2650.stack\[10\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07814_ _02188_ _02222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05925__B1 _05777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08794_ _02101_ _03044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_85_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_16_wb_clk_i_I clknet_4_4_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07745_ _02157_ _02164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05940__A3 _05793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10277__A2 _04412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11474__A1 _00740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11474__B2 _00519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07676_ _02091_ _02092_ _02098_ _02099_ _00034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_80_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09415_ _02730_ _02580_ _03598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06627_ as2650.holding_reg\[0\] _00654_ _01071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_13_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10029__A2 _04180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06558_ _00961_ _01002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_142_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_139_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09346_ _02143_ _02437_ _02147_ _03545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_139_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09277_ _03475_ _03491_ _03492_ _00242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_142_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06489_ _00932_ _00933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_103_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08228_ _02519_ _02531_ _02535_ _02540_ _00145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_33_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06653__B2 _01096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11700__CLK clknet_leaf_114_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_14_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08159_ _02488_ _02489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_180_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11201__I _01869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06405__A1 _00476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10201__A2 _00740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11170_ as2650.stack\[13\]\[2\] _05266_ _02002_ as2650.stack\[15\]\[2\] _05267_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_161_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10121_ as2650.addr_buff\[3\] _04124_ _04126_ _04202_ _04273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__06956__A2 _00655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_55_wb_clk_i_I clknet_4_12_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_5612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output68_I net68 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10052_ _04118_ _04120_ _04202_ _04206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_7_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_5634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11076__C _05174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06184__A3 _00547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05931__A3 _05779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11465__A1 _04620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10268__A2 _02964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10954_ net69 _05055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__07133__A2 _00962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10885_ _04199_ _04961_ _04897_ _04989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_31_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11217__A1 _05160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06892__A1 as2650.holding_reg\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09497__B _03660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09830__A1 _03987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07796__I _02206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11506_ _04948_ _04463_ _05555_ _00408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_156_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_94_wb_clk_i_I clknet_4_10_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11437_ _01721_ _05499_ _05504_ as2650.r123\[2\]\[0\] _05505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_144_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11111__I _05165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09433__I1 _03609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08397__A1 _02684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11368_ as2650.r123_2\[3\]\[6\] _05453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10319_ _04448_ _04449_ _04450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11299_ _02861_ _02810_ _05390_ _05391_ _00759_ _05392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_112_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08149__A1 as2650.stack\[8\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05860_ _05713_ _05714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_120_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09649__A1 _03793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09649__B2 _03811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11456__A1 _01622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07530_ as2650.stack\[7\]\[14\] _01959_ _01944_ as2650.stack\[6\]\[14\] _01960_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_35_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06875__I _01156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07461_ as2650.stack\[3\]\[11\] _01862_ _01863_ as2650.stack\[0\]\[11\] _01753_ as2650.stack\[1\]\[11\]
+ _01894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_50_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08872__A2 _03113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09200_ _03415_ _03419_ _03420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_06412_ _00824_ _00857_ _00609_ _00858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_17_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07392_ _01826_ _01827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11208__B2 as2650.stack\[3\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_148_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09131_ _03322_ _03353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06343_ _00792_ _00793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__09416__A4 _00768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09821__A1 _03978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08624__A2 _00769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09062_ _03189_ _03257_ _03287_ _03288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_147_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06635__A1 _01077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06274_ _00727_ _00728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_147_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_159_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_96_wb_clk_i clknet_4_9_0_wb_clk_i clknet_leaf_96_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_129_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_147_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08013_ _02109_ _02376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_116_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09424__I1 _03267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_190_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08388__A1 as2650.stack\[2\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06115__I _00524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10195__A1 _00753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10195__B2 _00473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07060__A1 _01341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09964_ _00961_ _04119_ _04120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07060__B2 _01498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08915_ _01303_ _03093_ _03159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08330__I _02626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09895_ _04049_ _04052_ _04053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__09888__A1 net62 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10498__A2 _05777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08846_ _03070_ _03093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08777_ _02473_ _03031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05989_ _00447_ _00448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_96_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07728_ _02143_ _02146_ _02147_ _02148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_72_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07115__A2 _01108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07659_ _02021_ _02084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08863__A2 _03098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06874__A1 _01306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10670__A2 _01814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10670_ as2650.stack\[9\]\[4\] _01814_ _01817_ as2650.stack\[8\]\[4\] as2650.stack\[10\]\[4\]
+ _01875_ _04780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_22_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_55_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09329_ _03037_ _03519_ _03531_ _03532_ _00254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_70_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_4_11_0_wb_clk_i_I clknet_3_5_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_194_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08615__A2 _01686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10958__B1 _05057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06626__A1 _01061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08505__I _02777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_193_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11222_ _03273_ _05125_ _05317_ _05318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_162_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_1686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_190_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11153_ _01219_ _05250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_150_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10104_ _04255_ _04103_ _04104_ _04256_ _01291_ _04257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_81_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11084_ _05176_ _05182_ _05183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_5420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09879__A1 _03987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10035_ _04181_ _04099_ _04190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_5464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10489__A2 _04589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_149_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06695__I _01120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11746__CLK clknet_leaf_113_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11986_ _00355_ clknet_leaf_77_wb_clk_i net67 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_186_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10110__A1 _03867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10937_ _04590_ _05030_ _05038_ _04891_ _05039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_72_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08854__A2 _03100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_189_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10868_ as2650.ivec\[4\] _04972_ _04841_ _04947_ _04873_ _04973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XPHY_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__11896__CLK clknet_leaf_96_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10799_ _04237_ _04894_ _04896_ _04905_ _04906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_129_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10413__A2 _04525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11610__A1 _00697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_157_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07290__A1 _01290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07042__A1 _01432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10680__I _04530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07593__A2 _02020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_3_6_0_wb_clk_i_I clknet_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06961_ _01058_ _01399_ _01400_ _01401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__11126__B1 _05223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08700_ _01999_ _02001_ _02143_ _02023_ _02971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_05912_ _05765_ _05766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_45_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09680_ _03796_ _01125_ _01126_ _03804_ _03805_ _03842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_4
X_06892_ as2650.holding_reg\[3\] _01167_ _01332_ _01333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_55_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08631_ _02902_ _02903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_27_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05843_ _05696_ _05685_ _05697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_95_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_82_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08562_ _01433_ _02835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_78_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07513_ _01824_ _01944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_35_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10101__A1 _04009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08493_ _00833_ _02741_ _02765_ _02584_ _02766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__08845__A2 _01010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10652__A2 _04748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07444_ as2650.stack\[15\]\[10\] _01874_ _01877_ as2650.stack\[14\]\[10\] _01878_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_149_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06320__A3 _00769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07375_ _01809_ _01810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09114_ _03300_ _03336_ _03337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_13_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06326_ _00753_ _00761_ _00776_ _00009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10404__A2 _04339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08325__I _02632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09270__A2 _03483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10076__B _04229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06257_ as2650.cycle\[3\] _00713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07281__A1 _00838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06084__A2 _00542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09045_ _01905_ _03273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_117_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10168__A1 _00556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06188_ _00542_ _00647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_102_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07033__A1 _01451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_176_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_191_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_85_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11619__C _00712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08781__A1 _02368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09947_ _03741_ _04104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_8_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08995__I _02086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09878_ _02611_ _01473_ _04036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_4026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11769__CLK clknet_leaf_92_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08829_ _00744_ _00937_ _03061_ _03076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_46_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10340__A1 _00737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06729__B _01135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10340__B2 _04465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11840_ _00223_ clknet_leaf_101_wb_clk_i as2650.stack\[7\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07404__I _01738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11771_ _00154_ clknet_leaf_91_wb_clk_i as2650.stack\[4\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_98 io_oeb[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_1945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10722_ as2650.stack\[11\]\[5\] _04822_ _01822_ as2650.stack\[10\]\[5\] _04831_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__10643__A2 _04749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10653_ _02852_ _05767_ _04763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_41_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05859__I _05712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07279__C _01007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10584_ _04688_ _04695_ _04696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_126_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09013__A2 _03067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10159__A1 _04077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_181_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07024__A1 _01433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11205_ as2650.stack\[2\]\[3\] _05296_ _05297_ as2650.stack\[0\]\[3\] _05301_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_123_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08772__A1 as2650.stack\[8\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11136_ _05221_ _05233_ _05234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_95_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11108__B1 _05205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10005__I _03661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_95_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11067_ as2650.stack\[2\]\[0\] _01940_ _01942_ as2650.stack\[0\]\[0\] _05165_ _05166_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XTAP_5261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_95_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07327__A2 _01740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08524__A1 as2650.stack\[11\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08524__B2 as2650.stack\[10\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10018_ as2650.addr_buff\[1\] _04173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_77_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_5294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10331__A1 _00826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_149_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11969_ _00338_ clknet_leaf_50_wb_clk_i net45 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_60_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06838__A1 _01263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10634__A2 _04702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06302__A3 _00585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_125_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07160_ _01597_ _01598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_105_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_160_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10398__A1 _02834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_121_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06111_ _00467_ _00569_ _00570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_9_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07263__A1 _01028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06066__A2 _00524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07091_ _01504_ _01529_ _01530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_51_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06042_ _00500_ _00494_ _00501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_133_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09004__A2 _03233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11347__B1 _01962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07015__A1 _05802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11347__C2 _01959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09801_ _02859_ _03872_ _03954_ _03960_ _00818_ _03951_ _03961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai222_1
XANTENNA__07566__A2 _01993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08763__A1 _02302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_99_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07993_ as2650.stack\[14\]\[0\] _02360_ _02201_ _02361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__10570__A1 as2650.stack\[7\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10570__B2 as2650.stack\[6\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09732_ _02856_ _03888_ _03892_ _03893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_140_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06944_ _01211_ _01373_ _01365_ _01354_ _01384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_112_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09704__I _02932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09712__B1 _03857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09712__C2 _03836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09663_ _02846_ _00683_ _03742_ _03819_ _03825_ _03826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_06875_ _01156_ _01316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10322__A1 _02903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08614_ _01422_ _01501_ _01589_ _02886_ _02887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_05826_ _05679_ _05680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_83_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09594_ _03726_ _00801_ _03756_ _03757_ _03758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__10873__A2 _04232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08545_ _00613_ _02818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_42_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10625__A2 _01839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08476_ _02745_ _00886_ _02598_ _02748_ _02749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_36_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09491__A2 _02546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08294__A3 _02602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07427_ _01854_ _01857_ _01860_ _01861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_123_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_40_wb_clk_i clknet_4_6_0_wb_clk_i clknet_leaf_40_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_91_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07358_ _01793_ _01794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09243__A2 _03443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07254__A1 _01257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06309_ _00759_ _00760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06057__A2 _00515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07289_ _01724_ _01725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_139_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07894__I _02059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09028_ _03258_ _03259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_139_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08004__B _02366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08754__A1 as2650.stack\[1\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06303__I _00606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06765__B1 _01206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10561__A1 _04671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08939__B _03115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output50_I net50 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08506__A1 _01770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10864__A2 _02758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_61_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11823_ _00206_ clknet_leaf_90_wb_clk_i as2650.stack\[8\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_73_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08809__A2 _03054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11274__C1 _01937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10616__A2 _04702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11754_ _00137_ clknet_leaf_81_wb_clk_i as2650.stack\[6\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09489__C _03655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10705_ _00978_ _04586_ _04105_ _04814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__10495__I _03745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07493__A1 _01920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11685_ _00068_ clknet_leaf_125_wb_clk_i as2650.stack\[10\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_186_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10636_ net58 net57 net56 net55 _04746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_167_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06048__A2 _00485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10567_ _04667_ _04678_ _04679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_154_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08993__A1 _03033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11934__CLK clknet_leaf_61_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10498_ net8 _05777_ _04611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_154_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08745__A1 _02394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07309__I _01744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06213__I _00608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11119_ as2650.stack\[1\]\[1\] _05153_ _05154_ as2650.stack\[3\]\[1\] _05217_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_46_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput6 io_in[34] net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_5080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10304__A1 _02332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11706__D _00089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06660_ _00939_ _01104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10855__A2 _04954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_52_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_188_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06591_ _00609_ _00947_ _01035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_36_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07979__I _02012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08330_ _02626_ _02636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10607__A2 _04702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09473__A2 _00687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08276__A3 _02550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06287__A2 _00681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07484__A1 _01735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08261_ _00602_ _02570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_177_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11280__A2 _02002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07212_ _01648_ _01649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_14_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08192_ _02506_ _02514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09225__A2 _03443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07236__A1 _01671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07143_ _01480_ _01487_ _01581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_173_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07787__A2 _01989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08984__A1 _03000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07074_ _05751_ _01360_ _01513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_146_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10791__A1 net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06025_ net72 as2650.cycle\[0\] _00484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_66_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05893__S1 _05713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07539__A2 _01959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08736__A1 as2650.stack\[1\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10543__A1 _02071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06211__A2 _00669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07663__B _02063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07976_ _01663_ _02345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_28_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10801__C _04554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09715_ _02607_ _03877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06927_ _01214_ _01353_ _01366_ _01368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_142_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11099__A2 _05190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09646_ _03794_ _03802_ _03808_ _03809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_99_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06858_ _01122_ _01299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_167_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09577_ _00638_ _00893_ _03741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_110_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06789_ _01065_ _01064_ _01210_ _01231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_97_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11807__CLK clknet_leaf_134_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08528_ as2650.stack\[13\]\[6\] _02785_ _02795_ as2650.stack\[12\]\[6\] _02801_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_42_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09464__A2 _02536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07475__A1 _01889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08672__B1 _01297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08459_ _02348_ _02732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__11271__A2 _05210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11470_ _04331_ _00950_ _05529_ _05530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_109_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09216__A2 _03428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11957__CLK clknet_leaf_20_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10421_ _04534_ _04535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08975__A1 _01658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09609__I net93 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_192_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10352_ _00725_ _01004_ _04474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_3_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10782__A1 _02952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05884__S1 _05736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10283_ _00941_ _01345_ _00515_ _04420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_4_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08727__A1 _02461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_183_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12022_ _00391_ clknet_leaf_38_wb_clk_i as2650.r123\[2\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_105_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10534__A1 _03876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06202__A2 _00660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09344__I _02650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10711__C _04819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10837__A2 _04940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07702__A2 _02062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_146_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07799__I _02200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11806_ _00189_ clknet_leaf_134_wb_clk_i as2650.stack\[15\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09455__A2 _03613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06269__A2 _00719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__11262__A2 _02814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11737_ _00120_ clknet_leaf_108_wb_clk_i as2650.stack\[0\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_124_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11114__I _01912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06208__I _00666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11668_ _00051_ clknet_leaf_128_wb_clk_i as2650.stack\[14\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_15_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11014__A2 _01131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10619_ as2650.stack\[6\]\[3\] _01781_ _01757_ as2650.stack\[4\]\[3\] _04730_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_89_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11599_ _03972_ _05636_ _05642_ _05643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_127_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08966__A1 _02932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07769__A2 _02172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10773__A1 _02115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06441__A2 _00516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10525__A1 _04630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09391__A1 as2650.stack\[6\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07830_ _02234_ _02190_ _02124_ _02235_ _02236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA__06878__I _01318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07761_ as2650.stack\[11\]\[5\] _02163_ _02176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_38_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05952__A1 _05745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05952__B2 _05708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09143__A1 as2650.r0\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09500_ _03665_ _03638_ _03666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06712_ as2650.addr_buff\[5\] _01155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_53_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07692_ as2650.stack\[13\]\[6\] _02062_ _02114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_38_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09694__A2 net93 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09431_ _03608_ _00280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06643_ _00460_ _00591_ _01087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_25_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09362_ _02076_ _03558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06574_ _01015_ _01017_ _01018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_36_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08313_ _02609_ _02620_ _02621_ _02622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_177_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09293_ _03033_ _03494_ _03503_ _03505_ _00245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_20_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_178_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08244_ _02552_ _00483_ _00729_ _02553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_192_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07209__A1 as2650.r0\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11005__A2 _00598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10863__I _01847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08175_ _02493_ _02501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_120_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05957__I _05789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_180_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08957__A1 _01597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07126_ as2650.r123\[1\]\[6\] _01116_ _01563_ _01207_ _01564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_146_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11556__A3 _00950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07057_ _01490_ _01495_ _01496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_47_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06983__A3 _00434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06008_ net72 _00467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09592__C _03755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10516__A1 _04626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09382__A1 _03571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10531__C _04643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07959_ _02236_ _02329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10103__I net41 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10970_ _03749_ _05058_ _05070_ _05071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_21_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09685__A2 _03845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09629_ _03730_ _03791_ _03792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_28_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07696__A1 _02116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08508__I _01736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output13_I net13 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__11244__A2 _05180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_145_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11522_ _00730_ _03639_ _05571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_141_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_84_wb_clk_i_I clknet_4_8_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11453_ _01932_ _05498_ _05513_ as2650.r123\[2\]\[5\] _05516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06671__A2 _01106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08948__A1 _01530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10404_ _03714_ _04339_ _04355_ _04518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__08243__I as2650.cycle\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11384_ as2650.stack\[9\]\[10\] _05464_ _05465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__10755__A1 _04400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_164_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10335_ _02850_ _04462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06423__A2 _00671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10266_ _02778_ _01024_ _03673_ _04405_ _00318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_84_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12005_ _00374_ clknet_leaf_52_wb_clk_i as2650.r123_2\[3\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08176__A2 _02497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09373__A1 _02110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06698__I net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06187__A1 _00645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10197_ _00548_ as2650.cycle\[12\] _04347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_39_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11180__A1 _05264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05934__A1 as2650.ins_reg\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_35_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09676__A2 net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_182_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08418__I _02693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07322__I _01757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09958__B _02894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_143_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08100__A2 _02430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06290_ _00739_ _00705_ _00741_ _00742_ _00011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_174_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06111__A1 _00467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_190_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08939__A1 _02933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10616__C _04333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10210__A3 _03649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09980_ _01607_ _04136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_89_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07992__I _02359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08931_ _03173_ _01422_ _03127_ _03174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_135_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08167__A2 _02495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09364__A1 _03231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08862_ _01102_ _01112_ _03108_ _03109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA_clkbuf_leaf_129_wb_clk_i_I clknet_4_0_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07813_ _02189_ _02220_ _02221_ _02210_ _00049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_29_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07914__A2 _02293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05925__A1 _05776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08793_ _03040_ _03041_ _03042_ _03043_ _00207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_96_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09116__A1 _00640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07744_ _02148_ _02163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_72_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12008__CLK clknet_leaf_117_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_183_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05940__A4 _05749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11474__A2 _02599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07675_ as2650.stack\[13\]\[4\] _02062_ _02063_ _02099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_25_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09414_ _03571_ _03589_ _03596_ _03597_ _00274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06626_ _01061_ _01067_ _01070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__11182__C _05278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09345_ _03543_ _03544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_90_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11226__A2 _01422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06557_ _00946_ _01001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_178_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08772__B _02481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09276_ _03214_ _03338_ _03340_ as2650.r123_2\[2\]\[7\] _03492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_193_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06488_ _00923_ _00924_ _00927_ _00931_ _00932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_138_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10985__A1 _00804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08227_ as2650.stack\[5\]\[11\] _02538_ _02540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07850__A1 _02053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_180_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_clkbuf_leaf_1_wb_clk_i_I clknet_4_1_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08158_ _02487_ _02488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_180_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07109_ _01544_ _01545_ _01546_ _01547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__06405__A2 _00843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08089_ _02329_ _02430_ _02431_ _02434_ _00112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__08998__I _02493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_162_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10120_ _04270_ _04271_ _04272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_122_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_164_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_192_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10051_ _04175_ _04178_ _04205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_114_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_27_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11162__A1 _05209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06311__I _00671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_180_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09107__A1 _03327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06184__A4 _00642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09622__I _00696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_166_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05931__A4 _05784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10768__I net63 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10953_ _05026_ _04700_ _05053_ _05054_ _00727_ _00356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_189_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10673__B1 _01755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10884_ _04987_ _04988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06341__A1 _00574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_185_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08094__A1 _02388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11505_ _04437_ _00751_ _05555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_157_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11436_ _05503_ _05504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_138_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09594__A1 _03726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08397__A2 _02681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11367_ _05452_ _00372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_158_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_153_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10318_ _03609_ _02903_ _04449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08701__I _02971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11298_ _01602_ _02960_ _02810_ _05391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_106_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_136_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_171_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08149__A2 _02477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09346__A1 _02143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10249_ _03165_ _04394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10171__C _04321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07317__I _01752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06221__I _00523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10900__A1 _04999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09649__A2 _03809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08321__A2 _02627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07460_ _01854_ _01891_ _01892_ _01893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_50_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10664__B1 _01751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08148__I _02473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06411_ _00833_ _00836_ _00854_ _00856_ _00857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_37_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11208__A2 _05302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06883__A2 _01303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07391_ _01825_ _01826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_31_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09130_ _03350_ _03351_ _03352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06342_ net3 _00792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08085__A1 _02325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_108_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09821__A2 _01428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10967__A1 _04802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09061_ _01953_ _03251_ _03278_ _03286_ _03287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_120_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06273_ _05678_ _00727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07832__A1 as2650.stack\[14\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_191_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_175_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08012_ _02091_ _02373_ _02374_ _02375_ _00094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_163_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10719__A1 _04540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_85_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10195__A2 _04340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11392__A1 as2650.stack\[9\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09963_ _04075_ _01692_ _04119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_103_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09337__A1 as2650.stack\[4\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08914_ _03147_ _03073_ _03157_ _03158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09894_ _04001_ _04000_ _04051_ _04052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_134_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07227__I _01663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08845_ _01120_ _01010_ _03092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_150_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06131__I _00589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07899__A1 as2650.stack\[10\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08776_ _02976_ _03029_ _03030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05970__I _05779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05988_ as2650.ins_reg\[3\] _00447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_26_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input12_I io_in[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09442__I _02529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07727_ _02022_ _02147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08058__I _02112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07658_ _02040_ _02083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_148_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06609_ _01033_ _01049_ _01052_ _01053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06874__A2 _01052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07589_ _00470_ _02016_ _02017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_159_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10258__I0 _04399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09328_ _03231_ _03523_ _03527_ _03532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08076__A1 _02318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10958__A1 _04814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10958__B2 _04794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11698__CLK clknet_leaf_123_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11080__B1 _01961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09259_ _03460_ _03471_ _03476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06626__A2 _01067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07823__A1 _01518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07823__B2 _02229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08007__B _02366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06306__I _00756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11221_ _00757_ _05294_ _05306_ _05316_ _05278_ _05317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_104_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10186__A2 _04325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09617__I _03654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11152_ _00842_ _05249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_49_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_161_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10272__B _03689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09328__A1 _03231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10103_ net41 _04256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_122_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11083_ _05177_ _05179_ _05181_ _05182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__11087__C _05185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11135__A1 _05222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10034_ _02205_ _04101_ _04188_ _04189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08000__A1 _02364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08677__B _02926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09352__I _02049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_99_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11985_ _00354_ clknet_leaf_77_wb_clk_i net66 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_95_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09500__A1 _03665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10936_ _04708_ _05033_ _05038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_16_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10110__A2 _04262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10867_ _04469_ _04972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_176_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_53_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10798_ _04610_ _04884_ _04903_ _04904_ _04905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_12_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07600__I _01729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_172_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07290__A2 _01725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11419_ as2650.stack\[9\]\[5\] _05478_ _05490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_193_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10177__A2 _04327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08431__I _02710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09319__A1 _02284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06960_ _01344_ _01398_ _01389_ _01400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__11126__A1 as2650.stack\[9\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input4_I io_in[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11126__B2 as2650.stack\[11\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05911_ _05764_ _05765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06891_ _05770_ _00664_ _01332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_132_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08630_ _02901_ _02902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_39_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06886__I _01077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05842_ _05688_ _05696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_39_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06553__A1 _00934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08561_ _01602_ _02834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__11429__A2 _03337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07512_ as2650.stack\[3\]\[13\] _01940_ _01941_ as2650.stack\[0\]\[13\] _01942_ as2650.stack\[1\]\[13\]
+ _01943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_08492_ _02764_ _02726_ _02727_ _02333_ _02765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
Xclkbuf_leaf_112_wb_clk_i clknet_4_3_0_wb_clk_i clknet_leaf_112_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07443_ _01876_ _01877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_165_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11840__CLK clknet_leaf_101_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06320__A4 _00770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07374_ _01737_ _01809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_149_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07510__I _01795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09113_ _03303_ _03335_ _03336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_148_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06325_ _00623_ _00499_ _00762_ _00771_ _00690_ _00775_ _00776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_109_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11062__B1 _05157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10404__A3 _04355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09044_ _03272_ _00229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_15_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06256_ _00711_ _00712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06126__I _00544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11990__CLK clknet_leaf_26_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_190_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07018__C1 _01456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06187_ _00645_ _05675_ _00646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__10168__A2 _00715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09437__I _02533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07033__A2 _01284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10707__A4 _04815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_172_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09881__B _03794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08781__A2 _03029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09946_ _00682_ _04103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_28_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09877_ _02611_ _01473_ _04035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_4027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09730__A1 _02854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08828_ _03057_ _03075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10312__S _04423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10340__A2 _02614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08759_ as2650.stack\[1\]\[6\] _03004_ _03016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11207__I _01863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11770_ _00153_ clknet_leaf_92_wb_clk_i as2650.stack\[4\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_99 io_oeb[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_109_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10721_ as2650.stack\[9\]\[5\] _01828_ _01825_ as2650.stack\[8\]\[5\] _04830_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_186_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10652_ _02619_ _04748_ _04761_ _04606_ _04762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_41_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_107_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07420__I _01788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10267__B _03692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10583_ _01776_ _04691_ _04694_ _04695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_155_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_139_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_194_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09549__A1 _00911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10159__A2 _04309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09347__I _03545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11204_ _05295_ _05299_ _05300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08772__A2 _03026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11135_ _05222_ _05232_ _05233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_122_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11108__A1 _01146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11108__B2 _03138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11066_ _05164_ _05165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_5251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_95_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_5262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_5273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10017_ _04169_ _04171_ _04172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_114_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08524__A2 _02782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10331__A2 _04457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11117__I _05158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10619__B1 _01757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08288__A1 _05696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09485__B1 _03649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11968_ _00337_ clknet_leaf_50_wb_clk_i net44 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_91_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10095__A1 _00719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_189_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10095__B2 _03995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10919_ _01904_ _04995_ _05007_ _03667_ _00882_ _05022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_177_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11899_ _00268_ clknet_leaf_72_wb_clk_i as2650.stack\[6\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08426__I _02705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07330__I _01765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08870__B _03115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11595__A1 _05638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06110_ _00568_ as2650.last_intr net75 _00569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_195_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07090_ _01505_ _01528_ _01529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_145_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07263__A2 _00427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08460__A1 _02732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06041_ _00453_ _00500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_86_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07486__B _01872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11347__A1 as2650.stack\[13\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08161__I _01988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08212__A1 _02527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09800_ _00688_ _03960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08763__A2 _02695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07992_ _02359_ _02360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_87_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10570__A2 _02799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06943_ _01375_ _01382_ _01383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09731_ _03887_ _03891_ _00533_ _03892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07933__C _02158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09712__A1 _02851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08515__A2 _01736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09662_ _03824_ _03810_ _03825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09712__B2 _03873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06874_ _01306_ _01052_ _01314_ _01315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_95_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10322__A2 _00795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07505__I _01830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08613_ _01097_ _01195_ _01249_ _01350_ _02886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_27_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05825_ as2650.ins_reg\[4\] _05679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_39_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09593_ _02745_ _00748_ _03757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_54_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08544_ _01462_ _02815_ _02817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08279__A1 _00660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10086__A1 _02212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11471__B _00518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08475_ _02746_ _02747_ _00598_ _00603_ _02748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_24_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07426_ as2650.stack\[7\]\[10\] _01858_ _01859_ as2650.stack\[5\]\[10\] _01860_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_23_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08336__I _02632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07357_ _01754_ _01793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10389__A2 _04504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11586__A1 _05413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06308_ _00758_ _00759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07254__A2 _01690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07288_ _01723_ _01724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_156_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_80_wb_clk_i clknet_4_10_0_wb_clk_i clknet_leaf_80_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_178_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09027_ _05677_ _03257_ _03246_ _03258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_191_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06239_ _00695_ _00696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_156_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_145_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11736__CLK clknet_leaf_108_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_1782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07006__A2 _01445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_1793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_191_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10010__A1 _04131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09951__A1 _02126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08754__A2 _03004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06765__A1 as2650.r123\[1\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09929_ _04074_ _04079_ _04080_ _04085_ _04086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_120_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_output43_I net43 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11510__A1 _01986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_189_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11822_ _00205_ clknet_leaf_112_wb_clk_i as2650.stack\[8\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09630__I _00538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11753_ _00136_ clknet_leaf_81_wb_clk_i as2650.stack\[6\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_42_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11274__B1 _01936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11274__C2 as2650.stack\[3\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10704_ _04808_ _04810_ _04812_ _04418_ _04813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_1787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08246__I _02554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08690__A1 _00951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11684_ _00067_ clknet_leaf_125_wb_clk_i as2650.stack\[10\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10635_ _02082_ _04701_ _04745_ _04645_ _00347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_126_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11577__A1 _02778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10566_ _04668_ _04648_ _04675_ _04677_ _00521_ _04678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_155_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10497_ _04608_ _04610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11329__A1 _05243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07402__C1 as2650.stack\[11\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08745__A2 _02996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10552__A2 _04659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11118_ _05215_ _05216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_1_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06771__A4 _01212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11049_ _05124_ _05148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_64_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput7 io_in[35] net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_5081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10304__A2 _04437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07325__I _01757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06590_ _00432_ _01034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_36_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12041__CLK clknet_leaf_9_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08260_ _02568_ _02569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08681__A1 _02951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08156__I _02470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07211_ as2650.r123\[0\]\[7\] as2650.r123_2\[0\]\[7\] _05709_ _01648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_144_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08191_ _02206_ _02513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_53_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07995__I _02359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07142_ _01575_ _01580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_9_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11759__CLK clknet_leaf_82_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07073_ _05764_ _01217_ _01512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08984__A2 _03222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_35_wb_clk_i_I clknet_4_6_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10791__A2 _05721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06024_ _00478_ _00482_ _00483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_160_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_160_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09933__A1 _03772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08736__A2 _02998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06747__A1 _00885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10543__A2 _04597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11466__B _02754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07975_ _00811_ net77 _02343_ _02344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_87_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06926_ _01214_ _01353_ _01366_ _01367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09714_ net89 _03876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_101_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09645_ _03797_ _03803_ _03807_ _00534_ _03808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_06857_ _01268_ _01255_ _01298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_28_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09576_ _03739_ _03740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06788_ _01227_ _01228_ _01229_ _01230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XTAP_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09449__B1 _03619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_184_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08527_ as2650.stack\[15\]\[6\] _02799_ _01745_ as2650.stack\[14\]\[6\] _02800_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_19_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08267__A4 _02575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08458_ _02730_ _02722_ _01037_ _00834_ _02731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_168_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08672__A1 _01141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08672__B2 _02853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07409_ _01775_ _01844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_clkbuf_leaf_74_wb_clk_i_I clknet_4_11_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08389_ _02678_ _02667_ _02671_ _02679_ _00167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__11559__A1 _02584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10420_ _00799_ _02570_ _04534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_136_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08424__A1 _02686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10231__A1 _00564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08975__A2 _03177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10351_ _00697_ _04470_ _04473_ _00335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_124_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08015__B _02356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10782__A2 _04097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10282_ _04418_ _04419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_2_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12021_ _00390_ clknet_leaf_35_wb_clk_i as2650.r123\[2\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_151_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08727__A2 _02712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06738__A1 _01173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10534__A2 _02055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09625__I _03724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_43_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11095__C _05192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05961__A2 _05734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10298__A1 _01262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11805_ _00188_ clknet_leaf_3_wb_clk_i as2650.stack\[15\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11247__B1 _05310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06269__A3 _00723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07466__A2 _01874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11736_ _00119_ clknet_leaf_108_wb_clk_i as2650.stack\[0\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08663__B2 _02932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11901__CLK clknet_leaf_73_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11667_ _00050_ clknet_leaf_132_wb_clk_i as2650.stack\[14\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08415__A1 as2650.stack\[1\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10618_ as2650.stack\[7\]\[3\] _01839_ _01752_ as2650.stack\[5\]\[3\] _04729_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_122_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11598_ _05413_ _05640_ _05635_ _05641_ _05642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_127_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10549_ _04077_ _03865_ _04660_ _04661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06977__A1 _00885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_170_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09915__A1 _00808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07764__B _02140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_119_wb_clk_i_I clknet_4_2_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10525__A2 _04637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09391__A2 _03577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09518__I1 _03672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07760_ _02091_ _02172_ _02173_ _02175_ _00042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_133_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05952__A2 _05761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06711_ _01132_ _01154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_38_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07691_ _02112_ _02113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07154__A1 _01316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09430_ as2650.ivec\[5\] _03285_ _03604_ _03608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06642_ _00593_ _01086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_129_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09361_ _03555_ _03544_ _03556_ _03557_ _00261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_52_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06573_ _01016_ _00977_ _01017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
Xclkbuf_leaf_19_wb_clk_i clknet_4_5_0_wb_clk_i clknet_leaf_19_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_61_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08312_ _02571_ _02621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_177_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08654__A1 _00843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09292_ as2650.stack\[2\]\[2\] _03504_ _03500_ _03505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_21_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08243_ as2650.cycle\[8\] _02552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_127_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10461__B2 _04332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_162_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07209__A2 _01542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08174_ _02488_ _02500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11005__A3 _05103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07125_ _01562_ _01563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_146_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_192_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_173_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11556__A4 _02735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06968__A1 _01180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10764__A2 _04845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07056_ _01413_ _01400_ _01495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_161_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09906__A1 _04045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06007_ _05728_ _00465_ _00466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_82_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_153_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06983__A4 _05770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09382__A2 _03562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07958_ _02327_ _02279_ _02328_ _02281_ _00087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_75_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06909_ _01096_ _01326_ _01349_ _01350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_99_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07889_ _02268_ _02280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_71_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09628_ _02054_ _03790_ _03791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__10320__S _04425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11924__CLK clknet_leaf_49_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09559_ _03722_ _03723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_62_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_164_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10452__A1 _03745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_180_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11521_ _02618_ _05566_ _05570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_141_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_169_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11452_ _01223_ _03473_ _05515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_184_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10204__A1 _03688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10403_ _02602_ _03712_ _03705_ _04516_ _04517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XANTENNA__08948__A2 _03177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09070__A1 _01980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11383_ _05455_ _05464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10755__A2 _00699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10334_ _02342_ _04457_ _04461_ _00330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_178_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06423__A3 _00768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07620__A2 _02045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10265_ _04404_ _04405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07076__S _05710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12004_ _00373_ clknet_leaf_120_wb_clk_i as2650.r123_2\[3\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_191_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09373__A2 _02653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10196_ _04339_ _04345_ _04346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_39_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06187__A2 _05675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_35_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_146_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10691__A1 _04794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11125__I _01761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06219__I _00529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07439__A2 _01858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10443__A1 _03722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11719_ _00102_ clknet_leaf_5_wb_clk_i as2650.stack\[12\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_187_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10994__A2 _05080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput10 io_in[7] net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_174_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09061__A1 _01953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09600__A3 _01018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_143_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_170_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08930_ _01429_ _03093_ _03172_ _03173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_135_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08861_ _03107_ _03108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07812_ as2650.stack\[14\]\[11\] _02208_ _02221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08792_ as2650.stack\[8\]\[4\] _03035_ _03031_ _03043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_57_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09116__A2 _03103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07743_ _02060_ _02161_ _02162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07674_ _02036_ _02097_ _02098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08875__A1 _01136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07513__I _01824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06625_ _01061_ _01062_ _01068_ _01069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_09413_ _02129_ _02514_ _03574_ _03597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__10682__A1 net60 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11035__I _05103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06556_ _00968_ _01000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09344_ _02650_ _03543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10434__A1 _04540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_181_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09275_ _03477_ _03486_ _03489_ _03490_ _03491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_166_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06487_ _00928_ _00930_ _00931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_107_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10985__A2 _05079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08226_ _02516_ _02531_ _02535_ _02539_ _00144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_148_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08344__I _02644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07850__A2 _02237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08157_ _02154_ _02485_ _02486_ _02487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_193_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07108_ _05780_ _05774_ _01516_ _01543_ _01546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_101_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08088_ as2650.stack\[0\]\[14\] _02419_ _02434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_134_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07039_ as2650.holding_reg\[5\] _01478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10315__S _04425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10050_ _04200_ _04201_ _04203_ _04204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_88_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_102_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_5669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_4946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_169_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07118__A1 _05732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10952_ as2650.ivec\[7\] _04972_ _04941_ _05028_ _04643_ _05054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_112_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10673__A1 as2650.stack\[13\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_186_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10673__B2 as2650.stack\[12\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10883_ _04929_ _04899_ _00893_ _04986_ _04987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_189_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10425__A1 _01786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10784__I _02772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05878__I _05731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10976__A2 _04701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11504_ _05553_ _04463_ _05554_ _00407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_89_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07841__A2 _02242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_185_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05852__A1 as2650.ins_reg\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11435_ _00640_ _01106_ _05502_ _05503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_156_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11366_ as2650.r123_2\[3\]\[5\] _05452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_158_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09594__A2 _00801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_152_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10317_ _05674_ _04399_ _04448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11297_ _05388_ _05389_ _05390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_98_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10248_ _03150_ _04387_ _04393_ _00312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_117_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10179_ net28 _00611_ _03646_ _03781_ _04330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_121_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10900__A2 _00809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08857__A1 _00695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09034__B _03263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10664__A1 as2650.stack\[6\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10664__B2 as2650.stack\[5\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06410_ _00511_ _00765_ _00855_ _00856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_07390_ _01755_ _01825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_97_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06341_ _00574_ _00788_ _00790_ _00791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_148_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07489__B _01872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08085__A2 _02430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09282__A1 as2650.stack\[2\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09060_ _03285_ _03252_ _03286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_124_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06272_ _00625_ _00717_ _00724_ _00726_ _00013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__08164__I _02493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08880__I1 _01127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08011_ _02174_ _02202_ _02366_ _02375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__05843__A1 _05696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09034__A1 _03261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_144_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07001__C _01052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_171_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09962_ _04026_ _04029_ _04117_ _04070_ _04118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA_fanout92_I net42 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08913_ _03074_ _03156_ _03157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_103_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09893_ _02106_ _02933_ _04050_ _04051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08844_ _01019_ _03073_ _03090_ _03091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_189_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07899__A2 _02274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05987_ _00445_ _00446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08775_ _02466_ _03029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_57_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_leaf_34_wb_clk_i clknet_4_7_0_wb_clk_i clknet_leaf_34_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_38_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07726_ _02145_ _02146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07657_ _02081_ _02082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_26_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07520__A1 _01766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06608_ _01051_ _01052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_129_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07588_ _00568_ as2650.last_intr net75 _02016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_107_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10407__A1 _00519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10258__I1 _04400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06539_ _00709_ _00642_ _00982_ _00983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_107_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09327_ as2650.stack\[4\]\[3\] _03521_ _03531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_159_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09273__A1 _03487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08076__A2 _02420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07399__B _01777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06087__A1 _00466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10958__A2 _05046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08074__I _02418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11080__A1 as2650.stack\[13\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09258_ _00835_ _03101_ _03475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_142_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11080__B2 as2650.stack\[12\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08209_ _02525_ _02522_ _02523_ _02526_ _00140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_09189_ _03377_ _03405_ _03409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_119_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_181_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11220_ _05264_ _05315_ _05316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08802__I _02121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07846__C _02047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10553__B _04664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07587__B2 _00579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11151_ _05242_ _05244_ _05247_ _05248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_194_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_output73_I net73 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07418__I as2650.r123\[0\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10102_ as2650.addr_buff\[3\] _04255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10272__C _03707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09328__A2 _03523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06322__I _00772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11082_ as2650.stack\[14\]\[0\] _05180_ _01962_ as2650.stack\[15\]\[0\] _05181_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_95_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07339__A1 _01770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08958__B _03122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11135__A2 _05232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10033_ _03824_ _04183_ _04187_ _04188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_133_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_5444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_5455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_5477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10894__A1 as2650.ivec\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10894__B2 _04975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06562__A2 _00634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08839__A1 _01277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08249__I _02557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11984_ _00353_ clknet_leaf_77_wb_clk_i net65 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_40_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09500__A2 _03638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10646__A1 _04454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10935_ _05036_ _04769_ _05037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_17_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10866_ _04790_ _04947_ _04970_ _04298_ _04971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_147_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_31_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__11642__CLK clknet_leaf_37_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10797_ _04331_ _04904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_158_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06078__A1 _00536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_121_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_157_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09016__A1 _03102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10019__I _04173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07290__A3 _01104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09808__I _03878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11792__CLK clknet_leaf_86_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11418_ _03561_ _05487_ _05488_ _05489_ _00386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_172_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07578__A1 _00817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10177__A3 _02811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11278__C _05159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11349_ _05437_ _05440_ _05441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_125_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11126__A2 _02142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08527__B1 _01745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05910_ as2650.r0\[3\] _05764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07772__B _02140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06890_ as2650.holding_reg\[3\] _00654_ _01330_ _01331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_67_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10885__A1 _04199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05841_ _05691_ _05694_ _05695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_12_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07750__A1 _02167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08560_ _00594_ _02833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08159__I _02488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07511_ _01791_ _01942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_63_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10637__A1 _03958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08491_ _00502_ _02764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_23_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07998__I _02187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07442_ _01875_ _01876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_126_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07373_ _01196_ _01808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_149_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09112_ _03305_ _03334_ _03335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06324_ _00774_ _00775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10357__C _03659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11062__A1 as2650.stack\[6\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07805__A2 _02208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11062__B2 as2650.stack\[4\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06407__I _00852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_191_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09043_ _03270_ as2650.r123_2\[0\]\[2\] _03271_ _03272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_164_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06255_ _00640_ _00711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09007__A1 _03239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07018__B1 _01453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06186_ _05669_ _00645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_128_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_150_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10168__A3 _03650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10573__B1 _02785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06142__I _00480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09945_ _00688_ _04102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08518__B1 _01756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09876_ _01609_ _01596_ _04034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_4006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_161_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09730__A2 _01303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08827_ _03072_ _03074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08758_ _02409_ _03011_ _03014_ _03015_ _00200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_2615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10628__A1 _01733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07709_ _02104_ _02129_ _01997_ _02130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_1903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08689_ _02960_ _01700_ _02961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__11665__CLK clknet_leaf_121_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_57_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10720_ _02779_ _04825_ _04828_ _04829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_92_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07701__I _02121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_158_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_161_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10651_ _05673_ _04755_ _04761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_35_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08018__B _02356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10582_ _01787_ _04692_ _04693_ _04694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_186_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08960__C _03127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10800__A1 _02571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06480__A1 _05714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09549__A2 _00574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08532__I _02777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10283__B _00515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11203_ as2650.stack\[6\]\[3\] _05296_ _05297_ as2650.stack\[4\]\[3\] _05298_ _05299_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_163_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11098__C _02819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06232__A1 _00498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11134_ _05228_ _05231_ _05232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11108__A2 _00789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11065_ _01771_ _01768_ _05164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_5230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05891__I _05718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_5252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10016_ _04170_ _04142_ _04171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_81_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06535__A2 _00978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10619__A1 as2650.stack\[6\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10619__B2 as2650.stack\[4\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11967_ _00336_ clknet_leaf_40_wb_clk_i net43 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09485__A1 _00465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08288__A2 _02335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09485__B2 _03651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10095__A2 _04245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11292__A1 net53 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10918_ _04584_ _05014_ _05020_ _05021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_32_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07611__I _02038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11898_ _00267_ clknet_leaf_72_wb_clk_i as2650.stack\[6\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_149_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09237__A1 _03174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10849_ _04588_ _04953_ _04954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_32_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11044__A1 _01277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08460__A2 _02727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06040_ _00490_ _00498_ _00499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_117_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08442__I _02710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11347__A2 _05178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_3_2_0_wb_clk_i clknet_0_wb_clk_i clknet_3_2_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_114_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07991_ _01999_ _02000_ _02272_ _02023_ _02359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_99_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07971__A1 _00938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09730_ _02854_ _01303_ _03890_ _03891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_141_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06942_ _01376_ _01377_ _01381_ _01382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_151_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10858__A1 _04226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09661_ _03743_ _03824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09712__A2 _03872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06873_ _01234_ _01307_ _01313_ _01051_ _01314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_132_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_94_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08920__B1 _03130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08612_ _02882_ _02884_ _02885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_23_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05824_ _05677_ _05678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_110_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09592_ _03728_ _03736_ _03754_ _03755_ _03756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_27_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08543_ _02815_ _01032_ _01454_ _02816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_54_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09476__A1 _03639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08279__A2 _00848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10086__A2 _03788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08617__I _02889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08474_ _00703_ _02747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_165_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_23_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_64_wb_clk_i_I clknet_4_14_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07425_ _01791_ _01859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_91_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11043__I _02764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07356_ as2650.stack\[14\]\[8\] _01746_ _01791_ as2650.stack\[13\]\[8\] _01792_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_164_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11586__A2 _04837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06307_ _00685_ _00758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07287_ _00477_ _00859_ _01723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_137_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09026_ _00838_ _03256_ _03257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06238_ _00510_ _00695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_156_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06169_ _00627_ _00628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_156_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09400__A1 _02087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10010__A2 _03976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09951__A2 _04101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09928_ _03894_ _04084_ _03761_ _04085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_120_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10323__S _04425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10849__A1 _04588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09859_ _04008_ _04017_ _04018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_8_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11510__A2 _05165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output36_I net36 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11821_ _00204_ clknet_leaf_112_wb_clk_i as2650.stack\[8\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_45_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09467__A1 as2650.stack\[5\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_164_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11274__A1 as2650.stack\[1\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11752_ _00135_ clknet_leaf_81_wb_clk_i as2650.stack\[6\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_14_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11274__B2 as2650.stack\[0\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07431__I _01824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06475__C _00920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_186_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10703_ _04811_ _04792_ _04812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11683_ _00066_ clknet_leaf_129_wb_clk_i as2650.stack\[12\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06047__I _00505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10634_ _04533_ _04702_ _04728_ _04743_ _04744_ _04745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_167_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11577__A2 _05621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10565_ _04226_ _04676_ _04677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_182_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09358__I _02066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06453__A1 _00500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08262__I _02570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10496_ _04608_ _04609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_170_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11329__A2 _02924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06205__A1 as2650.ins_reg\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07402__B1 _01827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_109_wb_clk_i_I clknet_4_3_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11117_ _05158_ _05215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_150_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07606__I _02033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11048_ _05128_ _05145_ _05146_ _05147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_5071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xinput8 io_in[5] net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_5082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_162_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11128__I _01816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_162_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09458__A1 as2650.stack\[5\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11291__C _03859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10312__I0 _04444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07341__I _01776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08681__A2 _02952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07210_ _05750_ _01515_ _01647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_18_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08190_ _02505_ _02508_ _02509_ _02512_ _00135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__09696__C _00551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10916__B _05018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07141_ _01059_ _01578_ _01579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_9_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06444__A1 _00822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10635__C _04645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07072_ _01357_ _01510_ _01511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_145_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06023_ _00479_ _00481_ _00482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_66_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_160_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08197__A1 as2650.stack\[6\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09933__A2 _04089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06747__A2 _00515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07974_ _02342_ _00630_ _02343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11466__C _02740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06420__I _00651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09713_ _00523_ _03827_ _03875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06925_ _01356_ _01365_ _01366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_95_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09644_ _03804_ _03805_ _03806_ _03807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_56_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06856_ _00437_ _01297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_132_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11482__B _03666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09575_ _01042_ _03739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_55_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09449__A1 _03550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06787_ as2650.holding_reg\[2\] _01228_ _01229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11256__A1 _04409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10059__A2 _01611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08526_ _02781_ _02799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08347__I _02135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08121__A1 as2650.stack\[0\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_180_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08457_ _00948_ _02730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_23_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08672__A2 _01034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11008__A1 _05102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07408_ _01837_ _01838_ _01842_ _01843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_184_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_167_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11703__CLK clknet_leaf_115_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08388_ as2650.stack\[2\]\[11\] _02676_ _02679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_11_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10826__B _04771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11559__A2 _02725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07339_ _01770_ _01774_ _01775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09621__A1 _03732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08424__A2 _02700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08082__I _02419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10231__A2 _00556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10350_ _04471_ _04472_ _00467_ _04473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_191_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09009_ as2650.stack\[7\]\[7\] _03228_ _03241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11853__CLK clknet_4_12_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10281_ _02772_ _04418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10519__B1 _01823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_191_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12020_ _00389_ clknet_leaf_105_wb_clk_i as2650.stack\[9\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08810__I _03056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07935__A1 _02161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07396__C1 _01830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10534__A3 _02038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_150_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10298__A2 _04432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08360__A1 _02519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_27_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11804_ _00187_ clknet_leaf_3_wb_clk_i as2650.stack\[15\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11247__A1 as2650.stack\[8\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11247__B2 as2650.stack\[11\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08257__I _00506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07161__I _01451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08112__A1 _02402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_11735_ _00118_ clknet_leaf_108_wb_clk_i as2650.stack\[0\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09860__A1 _02107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08663__A2 _01611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06674__A1 _00999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11666_ _00049_ clknet_leaf_121_wb_clk_i as2650.stack\[14\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_35_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10617_ _04583_ _04716_ _04718_ _04727_ _04728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__08415__A2 _02697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11597_ _05221_ _04696_ _05641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10222__A2 _04359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10548_ _03876_ _03866_ _04660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_170_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06977__A2 _00766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10479_ _00809_ _03821_ _04591_ _04592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_142_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08179__A1 _02327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09816__I net35 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09915__A2 _01693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07926__A1 as2650.stack\[11\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_170_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_97_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_111_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06240__I _00696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06710_ _01136_ _01137_ _01152_ _01153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_133_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07690_ _05682_ _02112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07154__A2 _01591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06641_ _01083_ _01084_ _01085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10697__I _00444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09360_ _02074_ _03548_ _03553_ _03557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06572_ as2650.addr_buff\[6\] _01016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_59_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08103__A1 as2650.stack\[0\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08311_ _02610_ _02614_ _02617_ _02619_ _02620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_127_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09291_ _03495_ _03504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09851__A1 _03870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08654__A2 _01090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_166_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08242_ _05698_ _00490_ _00614_ _02550_ _02551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_53_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_59_wb_clk_i clknet_4_15_0_wb_clk_i clknet_leaf_59_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_193_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08173_ _02323_ _02489_ _02494_ _02499_ _00131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__11876__CLK clknet_leaf_99_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09603__A1 _03766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08116__B _02446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11321__I _00756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07124_ _01533_ _01536_ _01561_ _01562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_101_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11410__A1 _02074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06415__I _00860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06968__A2 _01188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07055_ _01092_ _01493_ _01494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09726__I _01002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06006_ _05700_ _00462_ _00464_ _00465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_66_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08630__I _02901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07917__A1 as2650.stack\[10\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07957_ as2650.stack\[10\]\[13\] _02278_ _02328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_116_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06908_ _01327_ _01337_ _01340_ _01348_ _01349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__11477__A1 _04346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07888_ _02278_ _02279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08342__A1 _02527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09627_ net9 _03790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_83_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06839_ _01252_ _01157_ _01253_ _01281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_43_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11229__A1 _02724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09558_ _02037_ _03722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08077__I _02418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08509_ _02781_ _02782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_169_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09842__A1 _03933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09489_ _02566_ _01712_ _02761_ _03655_ _03656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_24_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11520_ _05556_ _05558_ _05568_ _03780_ _05569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_145_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09410__B _03574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11451_ _05512_ _05514_ _00394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_127_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10275__C _04405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06408__A1 _00848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10402_ _02551_ _02556_ _03702_ _04516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__11401__A1 as2650.stack\[9\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10204__A2 _03714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11382_ _02672_ _05457_ _05461_ _05463_ _00376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_194_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10333_ _00737_ _04460_ _04343_ _04458_ _04461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_124_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11387__B _05461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10264_ _00695_ _04404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_79_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07908__A1 _02174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11818__D _00201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12003_ _00372_ clknet_leaf_59_wb_clk_i as2650.r123_2\[3\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_133_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10195_ _00753_ _04340_ _04342_ _04344_ _00473_ _04345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_65_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06060__I _00518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08696__B _02894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11468__A1 _02578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11749__CLK clknet_leaf_88_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09371__I _02100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11406__I _05460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06895__A1 _01230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10691__A2 _04793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11899__CLK clknet_leaf_72_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09833__A1 _02612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11718_ _00101_ clknet_leaf_134_wb_clk_i as2650.stack\[12\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_147_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10466__B _04530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_147_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput11 io_in[8] net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_128_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11649_ _00032_ clknet_leaf_134_wb_clk_i as2650.stack\[13\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11141__I _00641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07072__A1 _01357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10980__I _05079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10913__C _04364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08450__I _02722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_174_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11156__B1 _03653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08860_ _03103_ _03107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_111_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_6_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07811_ _02219_ _02220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_57_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_106_wb_clk_i clknet_4_3_0_wb_clk_i clknet_leaf_106_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_135_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08791_ _02097_ _03029_ _03042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09116__A3 _03338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11459__A1 _05517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07742_ _02160_ _02161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09281__I _03495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_96_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10667__C1 as2650.stack\[2\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07673_ _02096_ _02097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08875__A2 _03111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09412_ as2650.stack\[6\]\[7\] _03585_ _03596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06624_ _01063_ _01064_ _01066_ _01067_ _01068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_129_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10682__A2 _04746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09343_ _01030_ _03542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06555_ _00998_ _00999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09824__A1 _03803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08627__A2 _01407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09274_ _03479_ _03483_ _03490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_146_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06486_ _00862_ _00929_ _00930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_166_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08225_ as2650.stack\[5\]\[10\] _02538_ _02539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_165_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_105_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10095__C _03777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08156_ _02470_ _02486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_174_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_162_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07107_ _05781_ _01516_ _01545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_146_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_31_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08087_ _02327_ _02430_ _02431_ _02433_ _00111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_106_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09456__I _02534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06810__A1 _00430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07038_ _00996_ _01458_ _01476_ _01477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_161_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_5604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11000__B _00679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_102_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08989_ _03028_ _03217_ _03224_ _03226_ _00220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_4925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07704__I net63 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08315__A1 _02610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10951_ _03662_ _05028_ _05051_ _05052_ _03832_ _05053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__10122__A1 _04270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06877__A1 _01016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05924__I0 as2650.r123\[1\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10882_ as2650.addr_buff\[0\] as2650.addr_buff\[1\] as2650.addr_buff\[2\] _04986_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_16_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06629__A1 _01068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08535__I _02807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11622__A1 net85 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11503_ _02860_ _00751_ _05554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_12_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05852__A2 _05705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11434_ _05697_ _05501_ _05502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__06055__I _05720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11365_ _05451_ _00371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_153_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_4_wb_clk_i clknet_4_1_0_wb_clk_i clknet_leaf_4_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__09366__I _02090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10733__C _04530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06801__A1 _01180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10316_ _04447_ _00326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11296_ _01599_ _02818_ _05134_ _02234_ _02812_ _05389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_10_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10305__I _04428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_191_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10247_ _04391_ _04392_ _04393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09346__A3 _02147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10178_ _02352_ _00899_ _04328_ _04329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_113_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08306__A1 _02341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10113__A1 _02218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10113__B2 _03830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11310__B1 _05269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10664__A2 _01780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_50_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10975__I _04404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_182_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09806__A1 _03951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10908__C _04752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06340_ _00781_ _00789_ _00474_ _00787_ _00790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XANTENNA__11613__A1 _05638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_175_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_148_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06271_ _00725_ _00690_ _00726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08010_ as2650.stack\[14\]\[4\] _02362_ _02374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_163_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05843__A2 _05685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_162_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07045__A1 _01478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10643__C _04752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08793__A1 _03040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07596__A2 _02001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09961_ _00792_ _01692_ _04117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11914__CLK clknet_leaf_73_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11129__B1 _05226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08912_ _01306_ _03075_ _03155_ _03156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_103_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09892_ _03957_ net12 _01464_ _02105_ _04050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout85_I net29 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08843_ _03074_ _03089_ _03090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_97_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10352__A1 _00725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06020__A2 _00462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08774_ _02050_ _03028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05986_ _00444_ _00445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_2_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07725_ _01991_ _02144_ _02145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_72_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10104__A1 _04255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10104__B2 _04256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06859__A1 _00437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10655__A2 _05761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07656_ _02080_ _02081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_53_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07520__A2 _01949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06607_ _01001_ _01050_ _01051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_74_wb_clk_i clknet_4_11_0_wb_clk_i clknet_leaf_74_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_94_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07587_ _00701_ _02009_ _02011_ _02014_ _00579_ _02015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_80_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10407__A2 _00893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10818__C _02334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09326_ _03033_ _03519_ _03529_ _03530_ _00253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_178_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06538_ _00956_ _00982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_22_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11604__A1 _05599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06087__A2 _00545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09257_ _03456_ _03474_ _00240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11080__A2 _05178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06469_ _00465_ _00913_ _00914_ _00915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_142_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_154_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08208_ as2650.stack\[6\]\[13\] _02517_ _02526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09188_ _03380_ _03404_ _03408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_193_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08139_ _02466_ _02475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_190_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08784__A1 _03033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_194_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11150_ net49 _05245_ _05246_ _05247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_122_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10591__A1 _02081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10101_ _04009_ _04247_ _04254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11081_ _01811_ _05180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_5401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output66_I net66 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10032_ _04186_ _00682_ _04104_ _04181_ _04105_ _04187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_114_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_102_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_5445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06562__A3 _00957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_99_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11983_ _00352_ clknet_leaf_77_wb_clk_i net64 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_4799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_95_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_4_4_0_wb_clk_i clknet_3_2_0_wb_clk_i clknet_4_4_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_10934_ _04395_ _03824_ _05036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_17_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09789__C _03948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10865_ _04948_ _04967_ _04969_ _02809_ _04970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__05889__I _05742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10796_ _03820_ _00689_ _04897_ _04902_ _04903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XPHY_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07275__A1 _05681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_160_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_15_wb_clk_i_I clknet_4_5_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11417_ as2650.stack\[9\]\[4\] _05476_ _05481_ _05489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_138_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07609__I net90 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07578__A2 _02005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06513__I _00956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11348_ _05209_ _05438_ _05439_ _05440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_181_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10582__A1 _01787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_180_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11279_ _05371_ _05372_ _05373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08527__A1 as2650.stack\[15\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08527__B2 as2650.stack\[14\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10334__A1 _02342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05840_ _05693_ _05694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__10885__A2 _04961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07344__I _01779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07510_ _01795_ _01941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_63_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08490_ _02756_ _02757_ _02762_ _02763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__10637__A2 _04746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07441_ _01779_ _01875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_126_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_54_wb_clk_i_I clknet_4_13_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07372_ as2650.r123\[0\]\[1\] _01807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__08175__I _02493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09111_ _03308_ _03333_ _03334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__07266__A1 _01664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06323_ _00773_ _00774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_160_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09042_ _03258_ _03271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_34_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_148_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06254_ _00694_ _00697_ _00708_ _00710_ _00002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_129_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09007__A2 _02495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_163_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07018__A1 _01432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07018__B2 _01299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06185_ _00625_ _00636_ _00643_ _00644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_117_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_121_wb_clk_i clknet_4_0_0_wb_clk_i clknet_leaf_121_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_116_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10573__A1 as2650.stack\[3\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09944_ _03751_ _04101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08518__A1 as2650.stack\[2\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08518__B2 as2650.stack\[0\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09875_ _02861_ _03850_ _04033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_189_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08826_ _03072_ _03073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_4029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10876__A2 _04979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_93_wb_clk_i_I clknet_4_8_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08757_ _02989_ _02695_ _02995_ _03015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_73_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05969_ _05773_ _00427_ _00428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_57_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07708_ _02128_ _02129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_2638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08688_ _02592_ _02960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_187_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10829__B _04819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07639_ net49 _02065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_13_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11651__D _00034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10650_ _04584_ _04753_ _04757_ _04759_ _04760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_179_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09309_ as2650.stack\[2\]\[7\] _03504_ _03493_ _03517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_10581_ as2650.stack\[15\]\[2\] _02908_ _02913_ as2650.stack\[13\]\[2\] _04693_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_194_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10800__A2 _02924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06480__A2 _05728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__11379__C _05461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07429__I _01795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08757__A1 _02989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11202_ _05159_ _05298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_120_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06333__I _00782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10564__A1 _01274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06232__A2 _00686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11133_ _05177_ _05229_ _05230_ _05231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_85_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_150_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11064_ _01941_ _05163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11395__B _05468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10015_ _02193_ _02940_ _04170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_5264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_5286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07164__I _01601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07732__A2 _01729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10619__A2 _01781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11966_ _00335_ clknet_leaf_69_wb_clk_i net72 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09485__A2 _03645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07496__A1 _01927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10917_ _03755_ _05016_ _05019_ _05020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__11292__A2 _05131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11897_ _00266_ clknet_leaf_96_wb_clk_i as2650.stack\[3\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_18_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_166_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10848_ _04175_ _04723_ _04616_ _04953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06508__I _00489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09237__A2 _03297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07248__A1 _01096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11044__A2 _02813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10779_ _03870_ _00699_ _04886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_121_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08996__A1 _03231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08723__I _02109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06471__A2 _00916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08748__A1 _02399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08748__B2 _03008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10555__A1 _02902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07990_ _02151_ _02222_ _02358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10921__C _04643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06941_ _05776_ _01380_ _01381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05982__A1 _05796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09173__A1 _05765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09660_ _03819_ _03820_ _03822_ _03823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06872_ _01309_ _01145_ _01027_ _01312_ _01313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__10858__A2 _04946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08920__A1 _01370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08611_ _00886_ _00461_ _02883_ _02884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_27_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08920__B2 as2650.r123_2\[1\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05823_ _05676_ _05677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09591_ _00799_ _03755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_36_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08542_ _02814_ _02815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_36_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10649__B _04725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09476__A2 _03640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08473_ _00952_ _02746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_78_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08119__B _02435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07424_ _01836_ _01858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_162_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06418__I _00863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09228__A2 _03446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07355_ _01790_ _01791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06306_ _00756_ _00757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_137_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07286_ _01717_ _01722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_148_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09025_ _03060_ _03063_ _03064_ _03066_ _03256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_136_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06237_ as2650.cycle\[4\] _00694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_163_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07249__I _01685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08739__A1 _03000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_1773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06168_ _00626_ _00627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_195_1784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10546__A1 _02851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09400__A2 _02514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06099_ as2650.cycle\[13\] net6 _00558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_120_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05992__I _00450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09927_ _04076_ _01696_ _04083_ _04084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_104_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11632__CLK clknet_leaf_36_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09858_ _03925_ _04011_ _04012_ _04016_ _04017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08911__A1 _03148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08809_ _01050_ _03054_ _03056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09789_ _02859_ _03894_ _03947_ _03948_ _03949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_3136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_185_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11820_ _00203_ clknet_leaf_113_wb_clk_i as2650.stack\[8\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09413__B _03574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11782__CLK clknet_leaf_88_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09467__A2 _03620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output29_I net29 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11751_ _00134_ clknet_leaf_88_wb_clk_i as2650.stack\[7\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_42_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11274__A2 _01934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_157_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10702_ _03750_ _04811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_41_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06328__I _00513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06150__A1 _00489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11682_ _00065_ clknet_leaf_129_wb_clk_i as2650.stack\[12\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_35_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10633_ _04529_ _04744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_122_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07868__B _02257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10564_ _01274_ _03744_ _04676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_139_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10785__A1 _04808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_194_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06453__A2 _00898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07650__A1 _02067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10495_ _03745_ _04608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07650__B2 _02075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07159__I _01569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06063__I _00521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06205__A2 _00447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_151_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11116_ _05209_ _05211_ _05213_ _05214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_111_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11047_ _00428_ _00680_ _02867_ _01139_ _00823_ _05146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_81_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08902__A1 _03110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_162_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput9 io_in[6] net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XTAP_5083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06913__B1 _01212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08718__I _02710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_52_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09458__A2 _03620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07622__I net79 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_146_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07469__A1 _01784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11949_ _00318_ clknet_4_6_0_wb_clk_i as2650.prefixed vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11144__I _00594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10312__I1 as2650.holding_reg\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06141__A1 _00508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08681__A3 _02335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08969__A1 _02836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_192_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07140_ _01576_ _01577_ _01578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__10916__C _04904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_173_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_145_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07071_ _01379_ _01510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06444__A2 _00858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06022_ _00480_ _00447_ _00481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_160_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10528__A1 _04620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_192_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09394__A1 _03550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07973_ _02341_ _02342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09146__A1 _03365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09712_ _02851_ _03872_ _03857_ _03873_ _00818_ _03836_ _03874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai222_1
X_06924_ _01361_ _01364_ _01365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_99_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09643_ _03804_ _03805_ _01002_ _03806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06855_ _01224_ _01296_ _00016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_55_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06755__I0 as2650.r123\[0\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09574_ _03723_ _05672_ _03738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_83_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06786_ _01067_ _01228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07532__I _01827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09449__A2 _03613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08525_ _02789_ _02796_ _02797_ _02798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_149_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11256__A2 _01458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08657__B1 _01142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11054__I _01855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08121__A2 _02445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10464__B1 _02758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08456_ _02725_ _02728_ _02729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_23_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09887__C _04004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07407_ _01765_ _01840_ _01841_ _01842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_149_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08387_ _02219_ _02678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_167_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07338_ _01768_ _01773_ net73 _01774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_149_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10767__A1 _02116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07632__A1 _02057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07269_ _01251_ _01693_ _01705_ _01293_ _01706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_10_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09008_ _03047_ _03233_ _03238_ _03240_ _00225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_151_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10280_ _04415_ _04416_ _04417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_156_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10519__A1 as2650.stack\[11\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10519__B2 as2650.stack\[10\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09385__A1 _02272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06199__A1 _00651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07396__B1 _01827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11192__A1 _01725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07935__A2 _02231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07396__C2 as2650.stack\[1\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07699__A1 _02113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07699__B2 _02120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06371__A1 as2650.addr_buff\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07442__I _01875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11803_ _00186_ clknet_leaf_16_wb_clk_i net54 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11247__A2 _01961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08648__B1 _01817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08112__A2 _02436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_11734_ _00117_ clknet_leaf_109_wb_clk_i as2650.stack\[0\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_186_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06674__A2 _01099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07871__A1 as2650.stack\[12\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11665_ _00048_ clknet_leaf_121_wb_clk_i as2650.stack\[14\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05897__I _05750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_174_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10616_ _04609_ _04702_ _04726_ _04333_ _04727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_15_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08273__I _00992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11596_ _05553_ _05637_ _05639_ _05640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__10758__A1 _00522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10547_ _04200_ _03960_ _04588_ _04659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_128_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_127_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06977__A3 _01416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10478_ _03787_ _03866_ _04591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08179__A2 _02500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09376__A1 as2650.stack\[3\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11183__A1 _03267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07617__I _02044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05937__A1 _05789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10930__A1 _05026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11583__B _05241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06640_ _01073_ _01084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_1604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07352__I _01787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06571_ _00429_ _01015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_1659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08639__B1 _01794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08103__A2 _02445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09300__A1 as2650.stack\[2\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08310_ _02618_ _02619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_55_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09290_ _02368_ _03502_ _03503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_61_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06114__A1 _00549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09851__A2 _02612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08654__A3 _00493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08241_ _00992_ _00747_ _02550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_60_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07862__A1 as2650.stack\[12\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09279__I _03493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08172_ as2650.stack\[7\]\[11\] _02497_ _02499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09603__A2 _03092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07123_ _01539_ _01560_ _01561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_118_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11410__A2 _05480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07054_ _01490_ _01492_ _01493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
Xclkbuf_leaf_99_wb_clk_i clknet_4_9_0_wb_clk_i clknet_leaf_99_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__10662__B _04770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07955__C _02281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06005_ _00463_ _00455_ _00464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__07378__B1 _01812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07917__A2 _02293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09119__A1 _03098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11049__I _05124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10921__A1 as2650.ivec\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10921__B2 _05002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07956_ _02230_ _02327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06907_ _01341_ _01343_ _01344_ _01347_ _01165_ _01348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_29_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07887_ _02277_ _02278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_56_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09626_ _00552_ _03789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06838_ _01263_ _01264_ _01014_ _01279_ _01280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__06353__A1 _00781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09557_ _03720_ _03721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11229__A2 _04786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06769_ _01210_ _01111_ _01211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_58_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08508_ _01736_ _02781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_180_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09488_ _00773_ _00785_ _03654_ _03655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_70_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09842__A2 _03935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10988__A1 _04439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08439_ as2650.stack\[15\]\[11\] _02714_ _02716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_145_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11820__CLK clknet_leaf_113_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11450_ _01449_ _05499_ _05513_ as2650.r123\[2\]\[4\] _05514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_156_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08093__I _02022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10401_ _04481_ _04514_ _04515_ _04506_ _00343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__06408__A2 _00850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11381_ as2650.stack\[9\]\[9\] _05462_ _05463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__11401__A2 _05476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_180_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10332_ _02847_ _04460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__11970__CLK clknet_leaf_39_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10263_ _00568_ _02606_ _04403_ _00317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_140_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_3_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11165__A1 _05216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12002_ _00371_ clknet_4_15_0_wb_clk_i as2650.r123_2\[3\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_78_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05919__A1 as2650.ins_reg\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10194_ _00778_ _02008_ _04343_ _04344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_87_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10912__A1 _04432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09652__I _03657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11468__A2 _04353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09530__A1 _00878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08333__A2 _02636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07172__I _01609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07541__B1 _01762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06895__A2 _01235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_56_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09601__B _03740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09833__A2 _03850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10979__A1 net71 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07844__A1 _02239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11717_ _00100_ clknet_leaf_134_wb_clk_i as2650.stack\[12\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_19_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11648_ _00031_ clknet_leaf_3_wb_clk_i as2650.stack\[13\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput12 io_in[9] net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_174_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11579_ _04652_ _02614_ _02965_ _05610_ _05624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_116_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_192_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11156__A1 _01150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11156__B2 _02851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08021__A1 _02381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10903__A1 _04709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07810_ _01363_ _02191_ _02192_ _02218_ _02219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_26_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08790_ _02473_ _03041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_61_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06583__A1 _01025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09562__I _02039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07741_ _02155_ _02160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_38_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11459__A2 _03491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09521__A1 _02552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10667__B1 _01817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_187_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10667__C2 _01875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07672_ _02094_ _02041_ _02095_ _02096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_168_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09411_ _03568_ _03589_ _03594_ _03595_ _00273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_77_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06623_ _00653_ _01067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_179_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09342_ _03050_ _03533_ _03540_ _03541_ _00258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_181_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06554_ _00921_ _00997_ _00998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_40_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08906__I _01310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10657__B _04763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09824__A2 _03982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08627__A3 _02876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09273_ _03487_ _03488_ _03489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07835__A1 as2650.stack\[13\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06485_ _00455_ _00929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_138_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08224_ _02529_ _02538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_165_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08155_ _02033_ _02485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_119_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_194_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11395__A1 _02686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07106_ _05774_ _01543_ _01544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08641__I _02784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08086_ as2650.stack\[0\]\[13\] _02427_ _02433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__10392__B _04501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07037_ _01154_ _01471_ _01475_ _00996_ _01476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_66_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06810__A2 _05808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11147__A1 _05243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_161_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08012__A1 _02091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_102_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06574__A1 _01015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08988_ _02364_ _03222_ _03225_ _03226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09472__I _03638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_180_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_4937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_99_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07939_ _02278_ _02315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_29_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10950_ _01926_ _04622_ _05033_ _03666_ _00882_ _05052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__06326__A1 _00753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09609_ net93 _03773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_16_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06877__A2 _00977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10881_ _04794_ _04976_ _04981_ _04984_ _04985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_16_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05924__I1 as2650.r123\[0\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08079__A1 _02321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09276__B1 _03340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08816__I _03062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07720__I _02139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07826__A1 _02222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_169_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11502_ _05681_ _05553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_40_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06336__I _00785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_156_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_172_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11433_ _01137_ _00954_ _05500_ _01292_ _05501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_103_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07876__B _02264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10189__A2 _00565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11364_ as2650.r123_2\[3\]\[4\] _05451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_137_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08551__I _02823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08251__A1 _00785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10315_ _04446_ _01478_ _04425_ _04447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_193_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06801__A2 _01188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11295_ _05243_ _02804_ _05387_ _05388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_152_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11138__A1 _03261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11138__B2 _05235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10246_ _04384_ _04392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08003__A1 _02368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10177_ net82 _04327_ _02811_ _04328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_78_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11866__CLK clknet_leaf_34_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09503__A1 _00901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08306__A2 _02336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06317__A1 _00766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10113__A2 _04111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11310__A1 as2650.stack\[10\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08857__A3 _03103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11310__B2 as2650.stack\[8\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09806__A2 _03867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11074__B1 _05172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11613__A2 _04440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11152__I _00842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06270_ as2650.cycle\[9\] _00725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06246__I _00544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_175_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_156_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08242__A1 _05698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08793__A2 _03041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07596__A3 _02003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09960_ as2650.addr_buff\[0\] _04116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_170_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11129__A1 as2650.stack\[10\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07077__I _01515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11129__B2 as2650.stack\[8\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08911_ _03148_ _03078_ _03154_ _03087_ _03155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_103_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09891_ _04047_ _04048_ _04049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_98_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09742__A1 _03886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08842_ _01100_ _03075_ _03088_ _03089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10352__A2 _01004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_83_wb_clk_i_I clknet_4_8_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08773_ _03020_ _03022_ _03023_ _03027_ _00203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_111_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05985_ _00443_ _00444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_85_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07724_ _01993_ _02144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_22_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10104__A2 _04103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11301__A1 _05801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06859__A2 _01252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07655_ net58 _02080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06606_ _00935_ _00939_ _01050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07586_ _01080_ _02013_ _02014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_41_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09325_ _02449_ _03523_ _03527_ _03530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_90_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06537_ _00973_ _00975_ _00980_ _00981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_126_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10407__A3 _00565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09256_ as2650.r123_2\[2\]\[5\] _03342_ _03473_ _03177_ _03474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_139_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06156__I _00614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_194_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06468_ _00774_ _00914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08481__A1 _02730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05914__S0 _05683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08207_ _02230_ _02525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_154_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09187_ _03145_ _03298_ _03407_ _00237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06399_ _00844_ _00845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_153_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09025__A3 _03064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10834__C _03780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11739__CLK clknet_leaf_113_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08138_ _02314_ _02468_ _02469_ _02474_ _00121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__07036__A2 _01474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08233__A1 as2650.stack\[5\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_146_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10040__A1 _02205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11011__B _00637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10040__B2 _03830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07587__A3 _02011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09981__A1 net88 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08784__A2 _03022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08069_ as2650.stack\[0\]\[8\] _02419_ _02421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_162_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06795__A1 _01233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10100_ _03789_ _04252_ _04145_ _04253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__10591__A2 _04646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11080_ as2650.stack\[13\]\[0\] _05178_ _01961_ as2650.stack\[12\]\[0\] _05179_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_89_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11889__CLK clknet_leaf_102_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10031_ _04173_ _04186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_5424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_102_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11540__A1 _02648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output59_I net86 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11982_ _00351_ clknet_leaf_76_wb_clk_i net63 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_90_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09930__I net37 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10933_ _04327_ _05030_ _05034_ _04606_ _05035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_44_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10864_ _04968_ _02758_ _04947_ _04534_ _04969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_108_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__11056__B1 _05154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10795_ _03824_ _04901_ _04902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_128_wb_clk_i_I clknet_4_0_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07275__A2 _05670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_184_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11416_ _03509_ _05480_ _05488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_172_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09972__A1 _04116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11347_ as2650.stack\[13\]\[7\] _05178_ _01962_ as2650.stack\[15\]\[7\] as2650.stack\[14\]\[7\]
+ _01959_ _05439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_180_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11278_ as2650.stack\[14\]\[5\] _01933_ _01936_ as2650.stack\[12\]\[5\] _05159_ _05372_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_79_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09724__A1 _00728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08527__A2 _02799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10229_ _04377_ _02333_ _04378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10334__A2 _04457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07625__I _02035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06553__A4 _00996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_23_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_clkbuf_leaf_0_wb_clk_i_I clknet_4_1_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12044__CLK clknet_4_4_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07440_ _01810_ _01874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_23_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10919__C _00882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06710__A1 _01136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11047__B1 _02867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07371_ _01709_ _01720_ _01806_ _00022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_149_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09110_ _03316_ _03332_ _03333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_149_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11598__A1 _05413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06322_ _00772_ _00773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_175_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07266__A2 _01137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08463__A1 _02731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09041_ _03145_ _03245_ _03248_ _03269_ _03270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_136_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06253_ _00709_ _00692_ _00710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_163_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_1922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07018__A2 _01011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08191__I _02206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06184_ _00639_ _00640_ _00547_ _00642_ _00643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XANTENNA__06704__I _00932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10022__A1 _04175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10573__A2 _02908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09943_ _04087_ _04099_ _03728_ _04100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_131_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08518__A2 _01745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09874_ _04025_ _03888_ _04031_ _04032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_100_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11485__C _00727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11522__A1 _00730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08825_ _00981_ _00983_ _03054_ _03072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_100_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11057__I _01940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05968_ _05790_ _00427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_08756_ as2650.stack\[1\]\[5\] _02998_ _03014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_72_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input10_I io_in[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07707_ _01980_ _02124_ _02127_ _02128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_2628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05899_ _05711_ _05753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__11932__D _00301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08687_ _02346_ _02902_ _02958_ _02959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_54_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07638_ _02051_ _01998_ _02061_ _02064_ _00031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_1938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06701__A1 _01143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07569_ _01996_ _01997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_41_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11589__A1 _02746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_167_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09308_ _02184_ _03502_ _03516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07257__A2 _01690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10580_ as2650.stack\[14\]\[2\] _04681_ _02914_ as2650.stack\[12\]\[2\] _04692_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_142_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10261__A1 _00795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09239_ _03435_ _03452_ _03457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07009__A2 _01422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08206__A1 _02521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10013__A1 _04167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11201_ _01869_ _05297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09954__A1 _02808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08757__A2 _02695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_181_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_194_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11132_ as2650.stack\[14\]\[1\] _05225_ _02002_ as2650.stack\[15\]\[1\] _05230_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06232__A3 _00689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09706__A1 _03836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_95_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11063_ _01870_ _05162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_5221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07445__I _01818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11513__A1 _01306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10014_ _04168_ _04169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_5254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_5265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07193__A1 _01555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11277__B1 _05310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11965_ _00334_ clknet_leaf_17_wb_clk_i as2650.alu_op\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10916_ _04610_ _05007_ _05018_ _04904_ _05019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_11896_ _00265_ clknet_leaf_96_wb_clk_i as2650.stack\[3\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_60_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11904__CLK clknet_leaf_72_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_189_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10847_ _04916_ _04947_ _04951_ _04326_ _04952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_158_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10778_ _00445_ _04884_ _03641_ _04885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_146_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10755__B _04105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10252__A1 _04394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_185_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08996__A2 _03222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10004__A1 _02195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10046__I _04199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10004__B2 _03968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08748__A2 _02996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06759__A1 _01135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10555__A2 _04649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_158_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11586__B _05624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06940_ _01379_ _01380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_141_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input2_I io_in[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05982__A2 _05801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07355__I _01790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10307__A2 _04440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06871_ _01310_ _00933_ _01144_ _01311_ _01312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_112_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08920__A2 _03163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08610_ _02872_ _02881_ _02883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05822_ _05675_ _05676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09590_ _03737_ _03738_ _03748_ _03753_ _03754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_82_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06931__A1 _00999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09570__I _03733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11268__B1 _05205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08541_ _01037_ _02814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_35_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08472_ _05681_ _02745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_110_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07423_ as2650.stack\[6\]\[10\] _01855_ _01856_ as2650.stack\[4\]\[10\] _01857_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_126_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07354_ _01789_ _01790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_71_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07958__C _02281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10243__A1 _04200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06305_ _00755_ _00756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_176_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07285_ _01099_ _01721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_137_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06998__A1 _05813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09024_ _03098_ _03245_ _03248_ _03254_ _03255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_164_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_163_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06236_ _00676_ _00580_ _00684_ _00693_ _00003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_156_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_1752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08739__A2 _03001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06167_ net3 _00626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10546__A2 _04587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_160_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_85_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06098_ _00466_ _00557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_85_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11927__D _00296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09926_ _04034_ _04037_ _04082_ _04083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_132_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09857_ _00629_ _04015_ _03817_ _04016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_100_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07175__A1 _01602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08808_ _00945_ _03054_ _03055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_150_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09788_ _00641_ _03948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_100_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08739_ _03000_ _03001_ _02701_ _03002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_2425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11750_ _00133_ clknet_leaf_113_wb_clk_i as2650.stack\[7\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10701_ _02952_ _04015_ _04809_ _04810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11681_ _00064_ clknet_leaf_129_wb_clk_i as2650.stack\[12\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_42_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06150__A2 _00594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08824__I _03070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10632_ _04620_ _04703_ _04741_ _04742_ _04640_ _04743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_122_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10234__A1 _04374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10563_ _04672_ _04674_ _04675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_155_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10785__A2 _04889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10494_ _04327_ _04592_ _04605_ _04606_ _04607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__07650__A2 _01998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09927__A1 _04076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07402__A2 _01830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11115_ as2650.stack\[6\]\[1\] _05212_ _05153_ as2650.stack\[5\]\[1\] _05213_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_150_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09155__A2 _03372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11046_ _00760_ _05143_ _05144_ _05145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_77_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_77_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08902__A2 _03145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_4372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08666__A1 _05695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11948_ _00317_ clknet_4_14_0_wb_clk_i as2650.last_intr vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_166_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06141__A2 _00599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11879_ _00248_ clknet_leaf_98_wb_clk_i as2650.stack\[2\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_20_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11017__A3 _05115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11160__I _01747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07070_ _01507_ _01374_ _01508_ _01509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_51_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_161_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06021_ _00463_ _00480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_103_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_195_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10528__A2 _04581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09394__A2 _03575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07972_ _00476_ _02341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_64_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09711_ _03744_ _03873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06923_ _01134_ _01219_ _01363_ _01020_ _01364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_136_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07157__A1 _01565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09642_ _03796_ _01118_ _01124_ _03805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
X_06854_ _01225_ _01295_ _01296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_151_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06904__A1 _00491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10700__A2 _00628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06785_ _05757_ _01227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_09573_ _00672_ _03737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_55_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08524_ as2650.stack\[11\]\[6\] _02782_ _01745_ as2650.stack\[10\]\[6\] _02797_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08657__A1 _01772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08657__B2 _01771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10464__A1 _03726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08455_ _02723_ _02726_ _02727_ _00883_ _02728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XANTENNA__10464__B2 _04553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07406_ as2650.stack\[14\]\[9\] _01781_ _01757_ as2650.stack\[12\]\[9\] _01841_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_168_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08386_ _02675_ _02667_ _02671_ _02677_ _00166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_51_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_177_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10216__A1 _04314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07337_ _01771_ _01772_ _01773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_195_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11559__A4 _02774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10767__A2 _04789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07268_ _01288_ _01704_ _01705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__06164__I _00622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09909__A1 _03837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06219_ _00529_ _00677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_3_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09007_ _03239_ _02495_ _03216_ _03240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07199_ _05765_ _01359_ _01510_ _05751_ _01636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_117_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10519__A2 _01835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09475__I _03641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06199__A2 _00657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07396__A1 as2650.stack\[2\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11192__A2 _04741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_132_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_82_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09909_ _03837_ _04065_ _04066_ _03786_ _00300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_120_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07148__A1 _01082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_output41_I net41 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08896__A1 _01286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07699__A2 _02092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07723__I _02142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11802_ _00185_ clknet_leaf_16_wb_clk_i net53 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06339__I _00451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08648__A1 as2650.stack\[14\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08648__B2 as2650.stack\[12\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10455__A1 _04428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10455__B2 _04568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_11733_ _00116_ clknet_leaf_111_wb_clk_i as2650.stack\[0\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06123__A2 _00580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11664_ _00047_ clknet_leaf_121_wb_clk_i as2650.stack\[14\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07871__A2 _02260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10207__A1 _03700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10615_ _04720_ _04722_ _04724_ _04725_ _04726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_167_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_4_3_0_wb_clk_i_I clknet_3_1_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11595_ _05638_ _04433_ _04435_ _05553_ _05639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_155_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06074__I _00532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10546_ _02851_ _04587_ _04658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_127_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10477_ _04376_ _04590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_6_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11029_ _00971_ _01097_ _05127_ _03781_ _05128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_110_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08887__A1 _01262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11340__C1 as2650.stack\[2\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07633__I _02059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10694__A1 _02094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06570_ _01013_ _01014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_92_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08639__A1 as2650.stack\[5\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08639__B2 as2650.stack\[4\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10446__A1 _02037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09300__A2 _03504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09851__A3 _03743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08654__A4 _00464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08240_ _00650_ _02546_ _02548_ _02549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_20_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10997__A2 _04701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08464__I _00950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07862__A2 _02258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08171_ _02321_ _02489_ _02494_ _02498_ _00130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_14_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_192_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07122_ _01540_ _01559_ _01560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_158_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_174_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10943__B _04395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07053_ _00500_ _01491_ _01410_ _01492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_175_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06004_ as2650.ins_reg\[2\] _00463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10662__C _04771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07808__I _02216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07378__B2 as2650.stack\[6\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07029__B _01035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09119__A2 _03298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06050__A1 _00502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_68_wb_clk_i clknet_4_9_0_wb_clk_i clknet_leaf_68_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07955_ _02325_ _02279_ _02326_ _02281_ _00086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_68_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06906_ _01081_ _01343_ _01346_ _01347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_68_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07886_ _02186_ _02137_ _02034_ _02277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_28_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09625_ _03724_ _03788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06837_ _01140_ _01276_ _01278_ _01279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_16_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06353__A2 _00801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_110_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09556_ _03719_ _03720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_43_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06768_ _05814_ _01210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_97_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10437__A1 _02906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08507_ _02779_ _02780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_70_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06699_ _01141_ _01142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09487_ _00879_ _02348_ _03654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_62_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08438_ _02675_ _02707_ _02711_ _02715_ _00180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_51_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09055__A1 _03174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08369_ _02196_ _02663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_71_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10400_ net23 _04480_ _04515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_137_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11380_ _05455_ _05462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06408__A3 _00853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07605__A2 _02020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10204__A4 _04353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06664__I0 as2650.r123\[0\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10070__C1 _00817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10331_ _00826_ _04457_ _04459_ _00329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_101_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07718__I _01988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10262_ as2650.last_intr _02606_ _04301_ _04403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_180_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11165__A2 _05260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12001_ _00370_ clknet_opt_2_0_wb_clk_i as2650.r123_2\[3\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_136_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10193_ _04341_ _04343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_78_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10912__A2 _05002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08869__A1 _00609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09530__A2 _00490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10676__B2 _01844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07541__A1 as2650.stack\[14\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07541__B2 as2650.stack\[13\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_34_wb_clk_i_I clknet_4_7_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06069__I net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_182_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11645__CLK clknet_leaf_32_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09294__A1 as2650.stack\[2\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11850__D _00010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_143_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11716_ _00099_ clknet_leaf_135_wb_clk_i as2650.stack\[12\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_124_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07844__A2 _02220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_175_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_187_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09046__A1 _01904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11647_ _00030_ clknet_leaf_2_wb_clk_i as2650.stack\[13\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_89_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11795__CLK clknet_leaf_123_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11578_ _01983_ _05611_ _05623_ _05076_ _00412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_156_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10600__A1 _03914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_170_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10529_ _04529_ _04642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11578__C _05076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06532__I as2650.addr_buff\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11156__A2 _02866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10903__A2 _05004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_73_wb_clk_i_I clknet_4_10_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_42_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06583__A2 _01026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07740_ _01984_ _02141_ _02150_ _02159_ _00038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_133_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08459__I _02348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07363__I _01777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09521__A2 _00547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10667__A1 as2650.stack\[1\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10667__B2 as2650.stack\[0\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07671_ _01927_ _02042_ _02095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09410_ _02119_ _02514_ _03574_ _03595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06622_ _01065_ _00989_ _01021_ _01066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_25_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_37_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06553_ _00934_ _00969_ _00984_ _00996_ _00997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_94_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09341_ _02129_ _02634_ _03518_ _03541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08088__A2 _02419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09285__A1 _02976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11092__A1 _00805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09272_ _01975_ _02234_ _03482_ _03488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__06707__I _00423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06484_ _00743_ _00928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_33_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_115_wb_clk_i clknet_4_2_0_wb_clk_i clknet_leaf_115_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__07835__A2 _02104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08223_ _02513_ _02531_ _02535_ _02537_ _00143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__07031__C _00944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_193_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08922__I _01436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08154_ _02329_ _02480_ _02481_ _02484_ _00127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_174_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11395__A2 _05467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07105_ _01542_ _01543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08085_ _02325_ _02430_ _02431_ _02432_ _00110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_106_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07036_ _01154_ _01474_ _01475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06271__A1 _00725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11147__A2 _04696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08012__A2 _02373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09753__I _02080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08987_ _02493_ _03225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06574__A2 _01017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_170_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_4938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07938_ _02196_ _02314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08369__I _02196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07273__I as2650.r123\[0\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10658__A1 _03960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_186_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07869_ _02251_ _02263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_29_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06326__A2 _00761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09608_ _03771_ _03772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_189_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10880_ _04916_ _04975_ _04983_ _03641_ _04984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_09539_ _00901_ _02004_ _03703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_71_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09276__A1 _03214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08079__A2 _02420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11083__A1 _05177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07826__A2 _02231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11501_ _05552_ _00406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_8_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_156_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10830__A1 _02619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_169_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_12_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11432_ _01013_ _00934_ _01055_ _05500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_7_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11363_ _05450_ _00370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08251__A2 _02549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_180_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_138_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06352__I _00800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10314_ _04428_ _04397_ _02609_ _04446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_113_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11294_ _05385_ _05386_ _02818_ _05134_ _05387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__11138__A2 _05189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10245_ _04255_ _04391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_140_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06014__A1 _00458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10176_ _04326_ _04327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_62_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11845__D _00005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10649__A1 _04394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09503__A2 _02555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06317__A2 _00767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08711__B1 _02977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11310__A2 _05180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07911__I _02277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11074__A1 as2650.stack\[9\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06527__I _00561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11074__B2 as2650.stack\[11\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10821__A1 _04725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08490__A2 _02757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_156_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07045__A3 _01483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08242__A2 _00490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07358__I _01793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06262__I _00551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06253__A1 _00709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07450__B1 _01882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07596__A4 _02023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11129__A2 _05225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08910_ _03149_ _03080_ _03153_ _03085_ _03154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_63_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09890_ net62 _01607_ _04048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_112_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10337__B1 _04457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08841_ _01032_ _03078_ _03086_ _03087_ _03088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__10888__A1 _04752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11810__CLK clknet_leaf_5_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08189__I _02511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08772_ as2650.stack\[8\]\[0\] _03026_ _02481_ _03027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05984_ _05703_ _00442_ _00443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_113_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07723_ _02142_ _02143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_26_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07654_ as2650.stack\[13\]\[3\] _02025_ _02079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10668__B _01786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11960__CLK clknet_4_7_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06605_ _01034_ _01036_ _01040_ _01048_ _01049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_53_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09258__A1 _00835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07585_ _00948_ _02012_ _00576_ _02013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_53_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09324_ as2650.stack\[4\]\[2\] _03521_ _03529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11065__A1 _01771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06536_ as2650.addr_buff\[7\] _00979_ _00980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_34_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06437__I _00849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09255_ _03459_ _03472_ _03473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_138_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06467_ _00694_ _00510_ _00913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__05914__S1 _05712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06492__A1 _00746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08206_ _02521_ _02522_ _02523_ _02524_ _00139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_09186_ as2650.r123_2\[2\]\[2\] _03342_ _03406_ _03163_ _03407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06398_ _00590_ _05702_ _00844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_120_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09025__A4 _03066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08137_ _02473_ _02474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08233__A2 _02538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06244__A1 _00492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10040__A2 _04111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_83_wb_clk_i clknet_4_8_0_wb_clk_i clknet_leaf_83_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_161_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08068_ _02419_ _02420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_150_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06795__A2 _01236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07019_ _01457_ _01458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_134_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09483__I _00973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10030_ _03789_ _04172_ _04184_ _04145_ _04185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_5414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06900__I _01086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09497__A1 _03662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11981_ _00350_ clknet_leaf_76_wb_clk_i net62 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_91_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10932_ _04604_ _05033_ _05034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08827__I _03072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07731__I _02044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10863_ _01847_ _04968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_92_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__11056__A1 as2650.stack\[5\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_38_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11056__B2 as2650.stack\[7\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10794_ _04899_ _04900_ _04901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_160_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_185_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_16_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06791__B _01232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08562__I _01433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06483__A1 _00558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11415_ _05460_ _05487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_103_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_177_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11346_ as2650.stack\[12\]\[7\] _02271_ _05438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_193_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11833__CLK clknet_leaf_27_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11277_ as2650.stack\[13\]\[5\] _05171_ _05310_ as2650.stack\[15\]\[5\] _05371_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_79_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10760__C _04819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10228_ _04376_ _00450_ _04377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_132_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07735__A1 _02154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08932__B1 _03130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10332__I _02847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10159_ _04077_ _04309_ _04310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_181_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11983__CLK clknet_leaf_77_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09488__A1 _00773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11295__A1 _05243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08737__I _02044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08160__A1 as2650.stack\[7\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07641__I _02066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06710__A2 _01137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11047__A1 _00428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07370_ _01721_ _01722_ _01719_ _01805_ _01806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__11047__B2 _01139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11598__A2 _05640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06321_ as2650.cycle\[5\] _00772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_149_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09660__A1 _03819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08463__A2 _02734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09568__I net93 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09040_ _03267_ _03262_ _03268_ _03269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06252_ as2650.cycle\[11\] _00709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06474__A1 _00556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08472__I _05681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06183_ _00641_ _00537_ _00631_ _00642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__10507__I _04534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09412__A1 as2650.stack\[6\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07423__B1 _01856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09963__A2 _01692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07974__A1 _02342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09942_ _03733_ _04099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout90_I net55 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09517__B _03677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07816__I net68 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09873_ _04026_ _04029_ _04030_ _04031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_135_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11522__A2 _03639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08824_ _03070_ _03071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_150_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_85_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08755_ _02405_ _03011_ _03012_ _03013_ _00199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_85_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05967_ _00423_ _00425_ _00426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_100_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11286__A1 _05189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07706_ _02126_ _02083_ _02127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08686_ _02954_ _02957_ _02351_ _02958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_26_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_130_wb_clk_i clknet_4_0_0_wb_clk_i clknet_leaf_130_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_54_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05898_ _05751_ _05752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07551__I _01664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07637_ as2650.stack\[13\]\[1\] _02062_ _02063_ _02064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_1928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11073__I _01819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06701__A2 _01025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06167__I net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07568_ _01985_ _01989_ _01995_ _01996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_39_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11706__CLK clknet_4_4_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09307_ _03047_ _03508_ _03514_ _03515_ _00249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_55_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11589__A2 _00951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06519_ _00872_ _00959_ _00962_ _00963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_166_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07499_ _01909_ _01910_ _01930_ _00026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09651__A1 _03789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09238_ _03189_ _03338_ _03456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10261__A2 _04388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09169_ _03366_ _03389_ _03390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_154_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_4_8_0_wb_clk_i_I clknet_3_4_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09403__A1 _03509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10417__I _04530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06217__A1 _05674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11200_ _01862_ _05296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_134_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11210__A1 _05300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09954__A2 _04008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11131_ as2650.stack\[13\]\[1\] _02142_ _05226_ as2650.stack\[12\]\[1\] _05229_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_output71_I net71 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09167__B1 _02223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09706__A2 _03867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11062_ as2650.stack\[6\]\[0\] _05156_ _05157_ as2650.stack\[4\]\[0\] _05160_ _05161_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XTAP_5211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_88_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10013_ _04167_ _04136_ _04168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_103_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_77_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_5255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10721__B1 _01825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_5288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11277__A1 as2650.stack\[13\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11964_ _00333_ clknet_leaf_17_wb_clk_i as2650.alu_op\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11277__B2 as2650.stack\[15\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10915_ _04391_ _04988_ _05017_ _05018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_2_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_32_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09890__A1 net62 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11895_ _00264_ clknet_leaf_96_wb_clk_i as2650.stack\[3\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_57_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11029__A1 _00971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10846_ _04949_ _04950_ _04806_ _04951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_73_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09642__A1 _03796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10777_ _04877_ _04884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_12_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06456__A1 _00720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09388__I _02506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10252__A2 _04387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_145_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07405__B1 _01752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06759__A2 _01021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11329_ _05243_ _02924_ _05418_ _05419_ _05420_ _05421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_64_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11586__C _05630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12011__CLK clknet_leaf_117_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07636__I _02046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_113_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11504__A2 _04463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06870_ _00439_ _00932_ _01311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07184__A2 _01589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08381__A1 as2650.stack\[2\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05821_ net5 _05675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_10_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_114_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06931__A2 _01351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11268__A1 _01463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08540_ _02812_ _02813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_94_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11268__B2 _02835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08669__C1 _02940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08467__I _00964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10315__I0 _04446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11729__CLK clknet_leaf_88_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08133__A1 _01991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08471_ _02737_ _02569_ _02739_ _02743_ _02744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_39_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_91_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07422_ _01795_ _01856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_165_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07353_ _01749_ _01789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_91_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08416__B _02694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09298__I _02096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06304_ _00754_ _00755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11440__A1 _01808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10243__A2 _04388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11440__B2 as2650.r123\[2\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07284_ _01719_ _01720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_148_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09023_ _01101_ _03251_ _03253_ _03254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06235_ as2650.cycle\[12\] _00692_ _00693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_1731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_145_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_191_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06166_ _00547_ _00625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_191_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06097_ _00555_ _00556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10951__B1 _05051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09925_ _01610_ _04081_ _04082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_131_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06450__I _00895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09856_ _04000_ _04014_ _04015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08807_ _03053_ _03054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_111_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09787_ _03763_ _03946_ _03947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_189_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06999_ _01433_ _01036_ _01437_ _01438_ _01439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_3127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11259__A1 _02610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08377__I _02670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08738_ _02688_ _03001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08124__A1 _02412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08669_ _02049_ _01141_ _01466_ _02100_ _02940_ _05682_ _02941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XTAP_1725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10700_ _02106_ _00628_ _04809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_109_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_42_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06686__A1 _00904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11680_ _00063_ clknet_leaf_131_wb_clk_i as2650.stack\[12\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10631_ _02758_ _04742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_139_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11531__I _02777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10234__A2 _00901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10562_ _00895_ _04673_ _04674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_126_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10493_ _04374_ _04606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_10_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_13_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09927__A2 _01696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08840__I _03056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11195__B1 _05288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07456__I _01351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06610__A1 _01013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11114_ _01912_ _05212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_123_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11045_ _02845_ _02842_ _05144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_5041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_162_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07166__A2 _00922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08363__A1 as2650.stack\[3\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_162_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10170__A1 _03677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11947_ _00316_ clknet_leaf_55_wb_clk_i as2650.addr_buff\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_33_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09863__A1 _03975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08666__A2 _00493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07469__A3 _01901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_189_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_178_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09620__B _03758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11878_ _00247_ clknet_leaf_99_wb_clk_i as2650.stack\[2\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_33_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10258__S _04385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10829_ _05673_ _04934_ _04819_ _04935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_32_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06429__A1 _00471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11422__A1 as2650.stack\[9\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09091__A2 _03313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_173_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06020_ _05699_ _00462_ _00479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_145_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_192_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_142_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06270__I as2650.cycle\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07971_ _00938_ _02339_ _02340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09710_ _03871_ _03872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06922_ _01362_ _01363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_136_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07157__A2 _01017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09581__I _01130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08354__A1 as2650.stack\[3\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09641_ _01041_ _03092_ _03804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_06853_ _01226_ _01249_ _01294_ _01295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_55_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10161__A1 _00546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06904__A2 _01091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09572_ _00795_ _03731_ _03735_ _03736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06784_ _00968_ _01226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_110_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08523_ as2650.stack\[9\]\[6\] _02785_ _02795_ as2650.stack\[8\]\[6\] _02796_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_64_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09854__A1 _03933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08657__A2 _01043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_184_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08454_ _00602_ _02727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_195_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06873__C _01051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07405_ as2650.stack\[15\]\[9\] _01839_ _01752_ as2650.stack\[13\]\[9\] _01840_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_162_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09606__A1 _03761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08385_ as2650.stack\[2\]\[10\] _02676_ _02677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_50_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09606__B2 _03769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08146__B _02474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_149_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11413__A1 _02087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07336_ _01742_ _01772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_109_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_176_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_176_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07093__A1 _00999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10621__C1 as2650.stack\[2\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07267_ _01133_ _01696_ _01703_ _01704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_136_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09006_ _02118_ _03239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06840__A1 _01016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06218_ _00472_ _00673_ _00676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08660__I _00792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_195_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07198_ as2650.r0\[3\] _01378_ _01635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_145_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11938__D _00307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06149_ _00607_ _00608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_2_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08593__A1 _00880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07396__A2 _01824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06180__I _00638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09908_ _04041_ _03720_ _04066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_154_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_134_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09839_ _03995_ _03997_ _03776_ _03998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_100_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_46_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10152__A1 _02549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output34_I net34 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11801_ _00184_ clknet_leaf_122_wb_clk_i as2650.stack\[15\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_55_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_162_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_3_1_0_wb_clk_i clknet_0_wb_clk_i clknet_3_1_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_2245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08648__A2 _01875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10455__A2 _04564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_11732_ _00115_ clknet_leaf_108_wb_clk_i as2650.stack\[0\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08835__I _03081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_2289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06123__A3 _00581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10586__B _04697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_11663_ _00046_ clknet_leaf_132_wb_clk_i as2650.stack\[14\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_41_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_126_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10614_ _03746_ _04725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11404__A1 as2650.stack\[9\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10207__A2 _03716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09073__A2 _03295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11594_ _02956_ _05638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10545_ _00446_ _04649_ _04653_ _04656_ _04657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_183_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10476_ _02846_ _04587_ _04588_ _04589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11848__D _00008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11210__B _05222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08584__A1 _02845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06090__I _00548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10391__A1 _03285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_63_wb_clk_i_I clknet_4_15_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11028_ _04409_ _01019_ _05126_ _00971_ _05127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_49_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10143__A1 net92 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11340__B1 _05223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11340__C2 _02387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10694__A2 _04704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09836__A1 _03793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08639__A2 _01790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10446__A2 _00513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11171__I _01811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08170_ as2650.stack\[7\]\[10\] _02497_ _02498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09064__A2 _03288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07121_ _01541_ _01552_ _01558_ _01559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_140_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08811__A2 _00927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07052_ _01420_ _01412_ _01491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_106_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11917__CLK clknet_leaf_73_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06003_ _00460_ _00461_ _00462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_161_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_192_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07378__A2 _01811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_142_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06050__A2 _00508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07954_ as2650.stack\[10\]\[12\] _02319_ _02326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07824__I _02230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06905_ _00884_ _01345_ _01346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_96_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10134__A1 _04004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07885_ _02044_ _02276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_68_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07535__C1 _01859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11477__A4 _05536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06889__A1 _01267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09624_ _02055_ _03787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06836_ _01277_ _01140_ _00944_ _01278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_55_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09555_ _03718_ _03719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_37_wb_clk_i clknet_4_6_0_wb_clk_i clknet_leaf_37_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_06767_ _01134_ _01200_ _01209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09827__A1 _03978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08506_ _01770_ _01774_ _02779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_09486_ _00502_ _00504_ _03653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__08655__I net74 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_108_wb_clk_i_I clknet_4_3_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06698_ net9 _01141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_145_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08437_ as2650.stack\[15\]\[10\] _02714_ _02715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_145_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11081__I _01811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08368_ _02527_ _02658_ _02659_ _02662_ _00163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_137_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07319_ _01754_ _01755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_149_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08299_ _02607_ _02608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_137_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10070__B1 _04211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06813__A1 _00430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10330_ _00737_ _02845_ _04343_ _04458_ _04459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__08390__I _02226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10070__C2 net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_30_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10261_ _00795_ _04388_ _04402_ _00316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07369__A2 _01800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08566__A1 _02833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12000_ _00369_ clknet_4_10_0_wb_clk_i as2650.r123_2\[3\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09763__B1 _03742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_132_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10192_ _00601_ _04341_ _04342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_156_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08318__A1 _01985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07734__I _02153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10125__A1 _04256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08869__A2 _03055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09530__A3 _00669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_41_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07541__A2 _01782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_55_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11715_ _00098_ clknet_leaf_135_wb_clk_i as2650.stack\[12\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_124_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11646_ _00029_ clknet_leaf_31_wb_clk_i as2650.r123\[0\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_35_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11577_ _02778_ _05621_ _05611_ _05622_ _05623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_168_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_10_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09396__I _03576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10600__A2 _03734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10528_ _04620_ _04581_ _04639_ _04640_ _04641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_122_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10335__I _02850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10459_ _03739_ _04571_ _04572_ _04225_ _04573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__08557__A1 _02807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10364__A1 _01101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12129_ net81 net13 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_123_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10116__A1 _04256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11313__B1 _05310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07670_ _02093_ _02094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_37_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10667__A2 _01814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06621_ _05734_ _01065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_92_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09809__A1 _03958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09809__B2 _03968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_20_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09340_ as2650.stack\[4\]\[7\] _03526_ _03540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06552_ _00970_ _00987_ _00995_ _00996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__11616__A1 _04460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09285__A2 _02681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08408__C _02694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06099__A2 net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09271_ _02346_ _03465_ _03487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06483_ _00558_ _00926_ _00927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__11092__A2 _00431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08222_ as2650.stack\[5\]\[9\] _02536_ _02537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_33_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08153_ as2650.stack\[8\]\[14\] _02467_ _02484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_147_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08424__B _02701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07104_ as2650.r123\[0\]\[6\] as2650.r123_2\[0\]\[6\] _05709_ _01542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_159_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07819__I _02226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08796__A1 as2650.stack\[8\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06723__I _01165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08084_ as2650.stack\[0\]\[12\] _02427_ _02432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_175_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10245__I _04255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07035_ _01473_ _01474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_164_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06271__A2 _00690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08548__A1 _01210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10355__A1 _00639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06023__A2 _00481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08986_ as2650.stack\[7\]\[1\] _03220_ _03224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_103_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07937_ _02161_ _02237_ _02313_ _02158_ _00081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_44_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07868_ _02220_ _02252_ _02257_ _02262_ _00063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_44_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08720__A1 _02456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06819_ _01254_ _01258_ _01260_ _01261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_09607_ _00538_ _00723_ _03771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_112_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07799_ _02200_ _02210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_37_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_186_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11607__A1 _05579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09538_ _00467_ _02016_ _03702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09276__A2 _03338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07287__A1 _00477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09469_ net26 _03636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_125_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11500_ as2650.r123\[3\]\[7\] _05552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_40_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10830__A2 _04921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11431_ _05498_ _05499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_12_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07729__I _02148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08334__B _02633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08787__A1 _02452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11362_ as2650.r123_2\[3\]\[3\] _05450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_193_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10594__A1 _02070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10313_ _04445_ _00325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_98_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11293_ net85 _02589_ _01724_ _05386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_106_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09944__I _03751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10244_ _01274_ _04387_ _04390_ _00311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_10_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06789__B _01210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06014__A2 _00472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10175_ _02608_ _04326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_154_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10649__A2 _00896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09503__A3 _03667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05913__S _05712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07514__A2 _01944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08711__A1 _02394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10758__C _03737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_186_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11762__CLK clknet_leaf_82_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07278__A1 _01103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11074__A2 _05171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_175_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_147_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10821__A2 _04925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11629_ net74 _05665_ _05668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_129_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08244__B _00729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07639__I net49 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08778__A1 as2650.stack\[8\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10585__A1 _04622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08242__A3 _00614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_183_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06253__A2 _00692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07450__A1 _01861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_87_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10337__A1 _04462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10337__B2 _00781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07202__A1 _01637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08840_ _03056_ _03087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_111_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10888__A2 _04979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08771_ _03025_ _03026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05983_ _05704_ _05693_ _00441_ _00442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XTAP_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07722_ _01782_ _02142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_61_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10949__B _04948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08702__A1 as2650.stack\[15\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07653_ _02077_ _02078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_25_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06604_ _01043_ _01045_ _01046_ _01047_ _01048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_187_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07584_ _00928_ _02012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_25_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09258__A2 _03101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08138__C _02474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09323_ _03028_ _03519_ _03525_ _03528_ _00252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06535_ _00976_ _00978_ _00979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08466__B1 _02738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11604__A4 _05646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09254_ _03460_ _03471_ _03472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_142_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10812__A2 _04917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06466_ _00911_ _00501_ _00703_ _00615_ _00912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_193_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08205_ as2650.stack\[6\]\[12\] _02517_ _02524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09185_ _03377_ _03405_ _03406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__06492__A2 _00469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06397_ _00837_ _00843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08154__B _02481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08136_ _02472_ _02473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_175_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10576__A1 _02780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_147_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_174_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06244__A2 _00457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08067_ _02418_ _02419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07993__B _02201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_150_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09764__I _00704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07018_ _01432_ _01011_ _01453_ _01299_ _01456_ _01426_ _01457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_150_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_172_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11635__CLK clknet_leaf_27_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_192_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_5415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10879__A2 _04982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08941__A1 _01460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_52_wb_clk_i clknet_4_13_0_wb_clk_i clknet_leaf_52_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_4714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_170_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08969_ _02836_ _03133_ _03208_ _03119_ _03209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_4736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11980_ _00349_ clknet_leaf_76_wb_clk_i net61 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_91_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09497__A2 _00623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10931_ _05031_ _05032_ _05033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_17_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08329__B _02633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10862_ _04879_ _04960_ _04964_ _04771_ _04966_ _04967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_147_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__11056__A2 _05153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10793_ _04847_ _04851_ _04898_ _04900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XPHY_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_34_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__10803__A2 _04878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__10594__B _02082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06791__C as2650.holding_reg\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06483__A2 _00926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07680__A1 as2650.stack\[13\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11414_ _03558_ _05473_ _05485_ _05486_ _00385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_138_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06363__I _00809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06235__A2 _00692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11345_ _05364_ _05435_ _05436_ _05437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_180_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09674__I net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_181_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_152_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11276_ _05365_ _05366_ _05369_ _05370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_180_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10227_ _03750_ _04376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07408__B _01842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08932__A1 _01387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10158_ _00631_ _00905_ _04309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_95_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10089_ as2650.addr_buff\[3\] _04242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_48_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09488__A2 _00785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11295__A2 _02804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10488__C _04432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08160__A2 _02488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06538__I _00956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11047__A2 _00680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06320_ _00763_ _00765_ _00769_ _00770_ _00771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XANTENNA__08999__A1 _02097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_175_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09660__A2 _03820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08463__A3 _02735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06251_ _00482_ _00545_ _00706_ _00707_ _00708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_148_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07671__A1 _01927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_121_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06273__I _05678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06182_ _00540_ _00530_ _00641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_129_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_1924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10558__A1 _01271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09412__A2 _03585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06226__A2 _00680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07423__A1 as2650.stack\[6\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11658__CLK clknet_leaf_124_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10951__C _03832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07974__A2 _00630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09941_ _04078_ _04097_ _04098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_132_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09872_ _04026_ _04029_ _03766_ _04030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_119_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08923__A1 _05813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08823_ _03066_ _03070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_97_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_161_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07037__C _00996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08754_ as2650.stack\[1\]\[4\] _03004_ _03005_ _03013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_85_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05966_ _00424_ _05785_ _00425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07705_ _02125_ _02126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_38_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08685_ _02951_ _02955_ _02956_ _02957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__11286__A2 _05363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05897_ _05750_ _05751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_38_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08151__A2 _02477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07636_ _02046_ _02063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06448__I _00893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_54_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07567_ _01994_ _01995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_41_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11038__A2 _05133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09100__A1 as2650.r0\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09306_ _03239_ _02673_ _03493_ _03515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_179_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06518_ _00478_ _00961_ _00962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_07498_ _01449_ _01911_ _01853_ _01929_ _01930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_139_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09651__A2 _03792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09237_ _03174_ _03297_ _03455_ _00239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_139_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06449_ _00894_ _00895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_142_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09168_ _05723_ _01380_ _03389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_135_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10549__A1 _04077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09403__A2 _03579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08119_ as2650.stack\[0\]\[5\] _02445_ _02435_ _02459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__11210__A2 _05305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09099_ _01544_ _03320_ _03321_ _01647_ _03322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_150_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09494__I _02807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11130_ _05224_ _05227_ _05228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_123_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09167__A1 _05724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09167__B2 _05743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11061_ _05159_ _05160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_5201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output64_I net88 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_5223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08914__A1 _03147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10012_ net87 _04167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XTAP_5234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_5245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_5256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10721__A1 as2650.stack\[9\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10721__B2 as2650.stack\[8\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_5289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08838__I _03077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07742__I _02160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11277__A2 _05171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11963_ _00332_ clknet_leaf_15_wb_clk_i as2650.alu_op\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_166_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10914_ _04242_ _04987_ _04570_ _05017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_75_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06153__A1 _00611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11894_ _00263_ clknet_leaf_95_wb_clk_i as2650.stack\[3\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_96_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11029__A2 _01097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10845_ _02195_ _04881_ _02204_ _04950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_144_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09669__I _03779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08573__I _01142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10776_ _04881_ _04882_ _04883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_13_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_157_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10788__A1 _04651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09642__A2 _01118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06456__A2 _00725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11800__CLK clknet_leaf_121_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_145_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06093__I _00551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_177_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07405__B2 as2650.stack\[13\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06759__A3 _01111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06821__I _01262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11328_ _02592_ _05242_ _05420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11950__CLK clknet_leaf_49_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05967__A1 _00423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10960__A1 _04811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11259_ _02610_ _05130_ _00847_ _05353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_140_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10712__A1 _04237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05820_ _05673_ _05674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08381__A2 _02673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06392__A1 _00476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07652__I _02076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11268__A2 _00789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08669__B1 _01466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08669__C2 _05682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10315__I1 _01478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08470_ _00763_ _02742_ _02743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__06144__A1 _00494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07421_ _01746_ _01855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_35_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07892__A1 _01984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07892__B2 _02282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09579__I _00681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07352_ _01787_ _01788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10779__A1 _03870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06303_ _00606_ _00754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11440__A2 _05499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07283_ _01718_ _01719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09022_ _01800_ _03252_ _03253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06234_ _00691_ _00692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_15_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10962__B _02331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09397__A1 as2650.stack\[6\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06165_ _00553_ _00621_ _00623_ _00624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_102_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_4_3_0_wb_clk_i clknet_3_1_0_wb_clk_i clknet_4_3_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_89_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_1765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_1787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05958__A1 _05808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06096_ _00554_ _00555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10951__A1 _03662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10951__B2 _05052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10253__I _02933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09924_ _01592_ _01594_ _01595_ _04081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_132_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07048__B _01483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_150_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09855_ _03957_ _01435_ _04013_ _04014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10703__A1 _04811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08806_ _00940_ _00651_ _03053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_41_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08658__I net85 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09786_ _03165_ _01445_ _03945_ _03946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_06998_ _05813_ _01147_ _01035_ _01438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_39_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05949_ _05798_ _05786_ _05803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_27_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08737_ _02044_ _03000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08124__A2 _02454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_167_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06178__I as2650.addr_buff\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08668_ _01608_ _02940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_1704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07619_ _02046_ _02047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_41_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08599_ net79 _01671_ _02872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_42_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05894__B1 _05747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10630_ _04731_ _04734_ _04740_ _01845_ _04741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_161_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_167_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_167_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08326__C _02633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10561_ _04671_ _04614_ _04669_ _04670_ _04673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_195_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10234__A3 _04375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_194_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10492_ _04604_ _04581_ _04605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10872__B _04676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__11195__A1 _03149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07737__I _02139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08342__B _02640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08060__A1 _02181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10942__A1 _04668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_53_wb_clk_i_I clknet_4_13_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11113_ as2650.stack\[4\]\[1\] _05210_ _05154_ as2650.stack\[7\]\[1\] _05211_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_146_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11044_ _01277_ _02813_ _05141_ _05142_ _05143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_110_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_5031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09560__A1 _00748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08363__A2 _02655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07472__I _01306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11946_ _00315_ clknet_leaf_54_wb_clk_i as2650.addr_buff\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07323__B1 _01758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09863__A2 _03976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07874__A1 _02231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11877_ _00246_ clknet_leaf_99_wb_clk_i as2650.stack\[2\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_33_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10828_ _04922_ _04934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_60_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10338__I _04464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06429__A2 _00870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11422__A2 _05476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10759_ _02351_ _04845_ _04867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_187_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_92_wb_clk_i_I clknet_4_8_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10630__B1 _04740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_145_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07929__A2 _02214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08051__A1 as2650.stack\[12\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10933__A1 _04327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11169__I _01782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_173_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07970_ _02332_ _00853_ _02338_ _02339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_142_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06921_ _01359_ _01362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08354__A2 _02653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06852_ _01251_ _01261_ _01289_ _01293_ _01294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_09640_ _03766_ _03803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_110_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06365__A1 _00550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_109_wb_clk_i clknet_4_3_0_wb_clk_i clknet_leaf_109_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__07382__I _01755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09571_ _03732_ _03734_ _03735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_49_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06783_ _01114_ _01225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_36_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09303__A1 as2650.stack\[2\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08522_ _02794_ _02795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09854__A2 _03963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08453_ _00879_ _00952_ _02726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_180_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_168_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07404_ _01738_ _01839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_168_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07331__B _01766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06726__I as2650.holding_reg\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08384_ _02665_ _02676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_36_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07335_ _01741_ _01771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__11413__A2 _05462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10621__B1 _01818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07093__A2 _01502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07266_ _01664_ _01137_ _01132_ _01702_ _01703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_137_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10621__C2 _01876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09005_ as2650.stack\[7\]\[6\] _03228_ _03238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06217_ _05674_ _00527_ _00624_ _00675_ _00004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_191_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07197_ _01632_ _01558_ _01633_ _01634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06840__A2 _00977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11177__A1 _05160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07557__I _01773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06148_ _00601_ _00517_ _00607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08042__A1 as2650.stack\[12\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_191_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11079__I _01877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08593__A2 _02865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06079_ _00537_ _00538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_120_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_78_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09907_ _04023_ _03788_ _04064_ _03977_ _04065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_63_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09542__A1 _00735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09838_ net35 _03996_ _03997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_150_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10152__A2 _02578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_189_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09769_ _03913_ _03929_ _03883_ _03930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_27_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11800_ _00183_ clknet_leaf_121_wb_clk_i as2650.stack\[15\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11101__A1 _02811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output27_I net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_2257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_11731_ _00114_ clknet_leaf_111_wb_clk_i as2650.stack\[0\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_155_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_187_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06636__I _00663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12001__CLK clknet_opt_2_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11662_ _00045_ clknet_leaf_126_wb_clk_i as2650.stack\[11\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_70_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10613_ _02855_ _04723_ _04724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11593_ _01675_ _01674_ _01685_ _05637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11404__A2 _05478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09947__I _03741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10544_ _04654_ _04655_ _04656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_122_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08281__A1 _00850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_182_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08820__A3 _03065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_104_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_170_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_157_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10475_ _03746_ _04588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07467__I _01815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08033__A1 _02276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11719__CLK clknet_leaf_5_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10915__A1 _04391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08584__A2 _02847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_7_wb_clk_i clknet_4_4_0_wb_clk_i clknet_leaf_7_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_155_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06595__A1 _00947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08800__B _03021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11869__CLK clknet_leaf_34_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11027_ _03794_ _01012_ _05126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09533__A1 _02585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08298__I _02012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06347__A1 _00611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07544__B1 _01973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11340__A1 as2650.stack\[1\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11340__B2 as2650.stack\[3\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09836__A2 _00723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11929_ _00298_ clknet_leaf_62_wb_clk_i net34 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_33_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_181_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10068__I net66 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07120_ _01553_ _01555_ _01557_ _01558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_70_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_118_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07051_ _01484_ _01489_ _01490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_173_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11401__B _05468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11159__A1 as2650.stack\[4\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06002_ _05772_ _00461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07377__I _01781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06281__I _00734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10906__A1 _04999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09772__A1 _02093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07953_ _02226_ _02325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09524__A1 _00616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06904_ _00491_ _01091_ _01345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__06338__A1 _00781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07884_ as2650.stack\[10\]\[0\] _02274_ _02275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10134__A2 _04285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07535__B1 _01856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07535__C2 as2650.stack\[1\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09623_ _03721_ _03784_ _03785_ _03786_ _00294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_95_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06835_ _01034_ _01277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_28_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06766_ _00999_ _01196_ _01208_ _00015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09554_ _03684_ _03698_ _03700_ _03717_ _03718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_24_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08505_ _02777_ _02778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_145_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06697_ _01039_ _01140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09485_ _00465_ _03645_ _03649_ _03651_ _03652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_93_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05849__B1 _05698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08436_ _02705_ _02714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06510__A1 _00947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_77_wb_clk_i clknet_4_11_0_wb_clk_i clknet_leaf_77_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_145_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08367_ as2650.stack\[3\]\[14\] _02645_ _02662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__11398__A1 _02151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07318_ net86 _01742_ _01754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_176_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08263__A1 _00645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_192_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08298_ _02012_ _02607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10070__A1 _04199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10070__B2 _00688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07249_ _01685_ _01686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__06813__A2 _05808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10260_ _00639_ _04392_ _04402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08015__A1 as2650.stack\[14\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09212__B1 _03431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_145_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09763__A1 _02855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08566__A2 _01700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09763__B2 _03886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10191_ _00734_ _00450_ _04341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_121_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11570__B2 _00839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09515__A1 _00865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__11322__A1 _05238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_98_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09530__A4 _02550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_28_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09451__B _03621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08846__I _03070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06794__C _01235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_182_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11714_ _00097_ clknet_leaf_127_wb_clk_i as2650.stack\[14\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06501__A1 _00744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_145_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11645_ _00028_ clknet_leaf_32_wb_clk_i as2650.r123\[0\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08581__I _02853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11576_ _04545_ _04552_ _05579_ _05622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_183_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10527_ _03915_ _04640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_155_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08006__A1 as2650.stack\[14\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10458_ _03739_ _04571_ _04572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_100_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_124_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08557__A2 _01498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09754__A1 _00881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10389_ _04481_ _04504_ _04505_ _04506_ _00340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__06568__A1 _00427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11561__A1 _00863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07925__I _02155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12128_ net81 net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_111_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11313__A1 as2650.stack\[13\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12047__CLK clknet_4_4_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11313__B2 as2650.stack\[15\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06620_ _00988_ _01064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_37_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06740__A1 _00592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06740__B2 _01082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_clkbuf_3_2_0_wb_clk_i_I clknet_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06551_ _00972_ _00975_ _00994_ _00995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_185_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11616__A2 _05575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09270_ _03479_ _03483_ _03486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06482_ _00529_ _00925_ _00926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_34_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08493__A1 _00833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06276__I _00729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08221_ _02529_ _02536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_147_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08152_ _02327_ _02480_ _02481_ _02483_ _00126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_140_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07048__A2 _01486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08245__A1 _00743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08491__I _00502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_158_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07103_ _05776_ _01514_ _01517_ _01541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_147_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10052__A1 _04118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08083_ _02423_ _02431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_134_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07034_ _01316_ _01453_ _01456_ _01319_ _01472_ _01473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_161_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08548__A2 _01135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09745__A1 _02080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11001__B1 _05099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06559__A1 _00714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_124_wb_clk_i clknet_4_0_0_wb_clk_i clknet_leaf_124_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__10355__A2 _04375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11552__A1 _03657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08440__B _02711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_102_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08985_ _03020_ _03217_ _03221_ _03223_ _00219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_130_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07936_ as2650.stack\[11\]\[14\] _02160_ _02313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_4929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11304__A1 _05209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07867_ as2650.stack\[12\]\[11\] _02260_ _02262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_28_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09606_ _03761_ _03764_ _03765_ _03768_ _03769_ _03770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_112_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08720__A2 _02712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06818_ _00423_ _01259_ _01260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_44_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07798_ as2650.stack\[14\]\[9\] _02208_ _02209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_44_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09537_ _02594_ _02602_ _03701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06749_ _01182_ _01191_ _01192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__11607__A2 _04444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09468_ _03571_ _03627_ _03634_ _03635_ _00290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08484__A1 _01143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10291__A1 _02332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08419_ as2650.stack\[1\]\[12\] _02697_ _02702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_169_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09399_ as2650.stack\[6\]\[3\] _03577_ _03587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_123_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11430_ _00514_ _00997_ _05498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_103_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08236__A1 _02527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10043__A1 _04181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_137_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09984__A1 _04001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11361_ _05449_ _00369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08787__A2 _02475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11240__B1 _02271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_180_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_192_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10594__A2 _04597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_180_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10312_ _04444_ as2650.holding_reg\[4\] _04423_ _04445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_152_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11292_ net53 _05131_ _05385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_152_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09736__A1 _03851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10243_ _04200_ _04388_ _04390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05974__B _00432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_175_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07745__I _02157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_191_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_26_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10174_ _03684_ _03715_ _04305_ _04324_ _04325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_154_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10104__C _01291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09503__A4 _03668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08711__A2 _02970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08576__I _02848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06722__A1 _01090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05930__C1 _05783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09267__A3 _03483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_182_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06096__I _00554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07278__A2 _01713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08475__A1 _02746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05908__S0 _05683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_54_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08227__A1 as2650.stack\[5\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11628_ _04444_ _05666_ _05667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10034__A1 _02205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08778__A2 _03026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10346__I _03692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11559_ _02584_ _02725_ _02728_ _02774_ _05605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_89_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08242__A4 _02550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10585__A2 _04696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_170_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10337__A2 _04463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11534__A1 _05561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07655__I net58 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05982_ _05796_ _05801_ _05804_ _00440_ _00441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_97_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08770_ _02388_ _02146_ _03024_ _03025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_84_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06961__A1 _01058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07721_ _02140_ _02141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_26_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08702__A2 _02972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08486__I _00784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07652_ _02076_ _02077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_130_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07390__I _01755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06603_ _00428_ _01044_ _01047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_80_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07583_ _00878_ _01080_ _05787_ _02010_ _02011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_20_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10030__B _04184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_168_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06534_ _00977_ _00978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_22_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09322_ as2650.stack\[4\]\[1\] _03526_ _03527_ _03528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__07269__A2 _01693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09663__B1 _03742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08466__B2 _00849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10273__A1 _03706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09253_ _03464_ _03470_ _03471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_146_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06465_ _00466_ _00911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_166_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08435__B _02711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_194_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08204_ _02511_ _02523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09184_ _03380_ _03404_ _03405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_147_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06396_ _00841_ _00842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_147_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10025__A1 _03794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09966__A1 _04116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08135_ _02153_ _01989_ _02471_ _02472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_159_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10025__B2 _03769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10256__I _02861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_193_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08066_ _01770_ _02249_ _02418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_190_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07017_ _01454_ _01455_ _01456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__09718__A1 _03876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07565__I _01992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11525__A1 _02625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_161_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_5416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_5438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08968_ _03078_ _03207_ _03208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_44_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06952__A1 as2650.holding_reg\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_102_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07919_ _02302_ _02297_ _02269_ _02303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_4759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_99_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08899_ _01249_ _03096_ _03144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_29_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07514__B _01866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10930_ _05026_ _05027_ _05032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_131_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_92_wb_clk_i clknet_4_8_0_wb_clk_i clknet_leaf_92_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_112_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10500__A2 _04612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_186_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10861_ _04752_ _04957_ _04965_ _04966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_71_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_92_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10792_ _04847_ _04851_ _04898_ _04899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_25_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08209__A1 _02525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06644__I _01087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07680__A2 _02025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09957__A1 _02126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11413_ _02087_ _05462_ _05481_ _05486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_172_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09957__B2 _02606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_193_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10567__A2 _04678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_opt_2_0_wb_clk_i_I clknet_4_10_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11344_ as2650.stack\[8\]\[7\] _05226_ _01962_ as2650.stack\[11\]\[7\] as2650.stack\[10\]\[7\]
+ _05180_ _05436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_138_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09709__A1 _03870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_180_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11275_ _05298_ _05367_ _05368_ _05369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__11516__A1 _03641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09185__A2 _03405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10226_ _00880_ _03650_ _01131_ _04375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_79_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07196__A1 _01541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08932__A2 _03163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10157_ _03685_ _04307_ _04308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07735__A3 _02034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10088_ _04068_ _04240_ _04241_ _00304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_48_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09623__C _03786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09488__A3 _03654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07499__A2 _01910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08696__A1 _02951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06755__S _05710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08448__A1 _02686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10255__A1 _04397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08999__A2 _03222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11460__I _02616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06250_ _00549_ _00707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_129_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06181_ _00510_ _00640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_8_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10558__A2 _05754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09865__I _02115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06226__A3 _00683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07423__A2 _01855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09940_ _04092_ _04096_ _04097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_104_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11507__A1 _00823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09871_ _03981_ _04027_ _04028_ _04029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08822_ _03065_ _03069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06934__A1 _05760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08753_ _02097_ _03001_ _03012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_61_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05965_ _05789_ _05790_ _05809_ _00424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_96_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07704_ net63 _02125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_26_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10679__C _04645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05896_ as2650.r0\[2\] _05750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08687__A1 _02346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08684_ _02597_ _02956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_94_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11286__A3 _05379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10494__A1 _04327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07635_ _02024_ _02062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07566_ _01991_ _01993_ _01994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_146_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09100__A2 _01542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09305_ as2650.stack\[2\]\[6\] _03496_ _03514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_55_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06517_ _00960_ as2650.idx_ctrl\[0\] _00961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_194_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07111__A1 _05758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07497_ _01890_ _01926_ _01928_ _01802_ _01929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_22_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09236_ as2650.r123_2\[2\]\[4\] _03340_ _03454_ _03107_ _03455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06448_ _00893_ _00894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_194_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09167_ _05724_ _01363_ _02223_ _05743_ _03388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06379_ _00491_ _00825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_108_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10549__A2 _03865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08118_ _02376_ _02442_ _02458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_174_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08611__A1 _00886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09098_ _05780_ _01543_ _01649_ as2650.r0\[0\] _03321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_135_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_194_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08049_ _02090_ _02405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_134_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05976__A2 _00434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09167__A2 _01363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11752__CLK clknet_leaf_81_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11060_ _05158_ _05159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_192_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07178__A1 _01598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10011_ _04068_ _04164_ _04166_ _00302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_5224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_5235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output57_I net89 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10721__A2 _01828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_185_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11962_ _00331_ clknet_leaf_20_wb_clk_i as2650.ins_reg\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08678__A1 _02926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10485__A1 _02057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10913_ _04604_ _05004_ _05015_ _04364_ _05016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_3888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11893_ _00262_ clknet_leaf_95_wb_clk_i as2650.stack\[3\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_60_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10844_ _02204_ net88 _04881_ _04949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_18_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07102__A1 _01520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10775_ _02125_ _04880_ _04802_ _04882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_40_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_158_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10788__A2 _04878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_82_wb_clk_i_I clknet_4_8_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08850__A1 _01097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06861__B1 _01298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07405__A2 _01839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11327_ _02951_ _00874_ _05135_ _05419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_141_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10960__A2 _05057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11258_ net52 _00873_ _05352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10209_ _03684_ _04358_ _04359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_39_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11189_ _05200_ _01350_ _05283_ _05284_ _03859_ _05285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_132_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10712__A2 _04817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08669__A1 _02049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08669__B2 _02100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10476__A1 _02846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06144__A2 _00602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07420_ _01788_ _01854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_78_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10228__A1 _04376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_162_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07351_ _01786_ _01787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_182_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10779__A2 _00699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06302_ _00662_ _00608_ _00585_ _00753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_07282_ _05677_ _01710_ _01717_ _01718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_149_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08841__A1 _01032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09021_ _03249_ _03252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_148_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06233_ _00553_ _00690_ _00691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__06217__C _00675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09595__I _00538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06164_ _00622_ _00623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11775__CLK clknet_leaf_92_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09397__A2 _03585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10400__A1 net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08432__C _02711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06095_ _00535_ as2650.cycle\[11\] _00554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_116_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05958__A2 _05770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06080__A1 _00529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10951__A2 _05028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09923_ _04078_ _03850_ _04080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_193_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_4_12_0_wb_clk_i_I clknet_3_6_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_127_wb_clk_i_I clknet_4_1_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09854_ _03933_ _03963_ _04013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_24_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06907__A1 _01341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09036__S _03259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10703__A2 _04792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08805_ _03050_ _03041_ _03051_ _03052_ _00210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09785_ _03943_ _03944_ _03945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06997_ _01436_ _01045_ _01437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_100_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08736_ as2650.stack\[1\]\[0\] _02998_ _02999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_73_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05948_ _05799_ _05802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_100_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10467__A1 _03726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08667_ _05687_ _00792_ _01042_ _01030_ _02076_ _02854_ _02939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_27_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05879_ _05732_ _05733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06135__A2 _00593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07618_ _01996_ _02046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06686__A3 _01128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08598_ _02805_ _02864_ _02870_ _02871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_41_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05894__A1 _05745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07549_ _01958_ _01910_ _01978_ _00028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__05894__B2 _05739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_195_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10560_ _04669_ _04670_ _04671_ _04614_ _04672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__08832__A1 _01143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_155_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09219_ _03420_ _03421_ _03438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_108_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10491_ _02824_ _04604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_10_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_178_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11195__A2 _02833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_123_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08060__A2 _02258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05949__A2 _05786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10942__A2 _05037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11112_ _01914_ _05210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_122_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_5010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11043_ _02764_ _05142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09454__B _03621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08899__A1 _01249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08849__I _03065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07753__I _02086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_5054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09560__A2 _02866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07166__A4 _00974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06374__A2 _00745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_4364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_4375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11945_ _00314_ clknet_leaf_54_wb_clk_i as2650.addr_buff\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09901__C _03925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07323__A1 as2650.stack\[5\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11648__CLK clknet_leaf_3_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07874__A2 _02263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11876_ _00245_ clknet_leaf_99_wb_clk_i as2650.stack\[2\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_3_7_0_wb_clk_i_I clknet_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10827_ _04668_ _04915_ _04932_ _04933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_32_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11798__CLK clknet_leaf_120_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10758_ _00522_ _04854_ _04865_ _03737_ _04866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__06429__A3 _00874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10630__B2 _01845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10689_ _04796_ _04797_ _04586_ _04798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_139_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08051__A2 _02390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10933__A2 _05030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06920_ _01357_ _05775_ _01218_ _01360_ _01361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_68_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09000__A1 as2650.stack\[7\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06851_ _01292_ _01293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09551__A2 _03712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06365__A2 _00713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11185__I _00696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09570_ _03733_ _03734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_55_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06782_ as2650.r123\[1\]\[2\] _01116_ _01222_ _01223_ _01224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_110_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09303__A2 _03504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08521_ _01754_ _02794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_82_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11110__A2 _05207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08452_ _02723_ _00870_ _02724_ _02725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_91_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07865__A2 _02260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05911__I _05764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07403_ as2650.stack\[10\]\[9\] _01812_ _01788_ _01838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_127_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09067__A1 _03202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08383_ _02213_ _02675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10529__I _04529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07334_ _01736_ _01769_ _01770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_91_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08814__A1 _00955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06825__B1 _05768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07265_ _01462_ _01040_ _01699_ _01701_ _00943_ _01702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_104_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10621__B2 as2650.stack\[0\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07838__I _02035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09004_ _03044_ _03233_ _03236_ _03237_ _00224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06742__I _01072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06216_ _00462_ _00644_ _00646_ _00674_ _00675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_07196_ _01541_ _01552_ _01633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10264__I _00695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06147_ _00605_ _00606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_145_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08042__A2 _02390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06078_ _00536_ as2650.cycle\[3\] _00537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06898__B _01058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09906_ _04045_ _04054_ _04061_ _04063_ _04064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_43_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_99_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_150_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07573__I _02000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09837_ net34 _03953_ _03996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__09542__A2 _00729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07553__A1 _01707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_115_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10152__A3 _03696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_150_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06189__I _00494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11028__C _00971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09768_ _03914_ _03725_ _03916_ _03928_ _03929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_46_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08719_ as2650.stack\[15\]\[4\] _02972_ _02986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_167_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09699_ _02070_ _01271_ _03861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_27_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11101__A2 _00760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08618__B _02890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_11730_ _00113_ clknet_leaf_109_wb_clk_i as2650.stack\[0\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__11940__CLK clknet_leaf_56_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05821__I net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10860__A1 _04326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_186_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11661_ _00044_ clknet_leaf_1_wb_clk_i as2650.stack\[11\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_148_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10612_ _00894_ _04723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08805__A1 _03050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_180_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11592_ net49 _05635_ _05636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__10883__B _00893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10543_ _02071_ _04597_ _04655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08820__A4 _03066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06292__A1 _00743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10474_ _04586_ _04587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08033__A2 _02392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09781__A2 _03940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08584__A3 _02851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_194_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06595__A2 _01038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07792__A1 _02189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08579__I net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10679__A1 _02094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11026_ _05124_ _05125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09533__A2 _02578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06347__A2 _00644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11340__A2 _05257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12041__D _00410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06827__I _01268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11928_ _00297_ clknet_leaf_63_wb_clk_i net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_33_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10851__A1 _04167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11859_ _00228_ clknet_leaf_31_wb_clk_i as2650.r123_2\[0\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_162_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_140_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10603__A1 _04391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07050_ _01485_ _01488_ _01489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_12_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_173_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06001_ _05771_ _00460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__11159__A2 _05210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_103_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09221__A1 _01569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06035__A1 _00492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09772__A2 net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_47_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11813__CLK clknet_leaf_111_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07952_ _02323_ _02315_ _02324_ _02317_ _00085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_151_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05906__I _05759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06903_ _01342_ _01333_ _01344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09524__A2 _02593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07883_ _02273_ _02274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_68_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06338__A2 _00783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07535__A1 as2650.stack\[3\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09622_ _00696_ _03786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06834_ _01269_ _01036_ _01270_ _01275_ _01276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_68_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06938__S net51 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11963__CLK clknet_leaf_15_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09553_ _03701_ _03706_ _03715_ _03716_ _03717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_06765_ as2650.r123\[1\]\[1\] _01197_ _01206_ _01207_ _01208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__09288__A1 _03028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08438__B _02711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08504_ _00865_ _02777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_149_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07342__B _01777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11095__A1 _02027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09484_ _02732_ _03650_ _03651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06696_ _01138_ _01139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05849__A1 _05681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_93_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05849__B2 _05702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08435_ _02672_ _02707_ _02711_ _02713_ _00179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_23_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06510__A2 _00953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08366_ _02525_ _02658_ _02659_ _02661_ _00162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_108_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11398__A2 _05467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07317_ _01752_ _01753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_123_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08297_ _00749_ _02606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08263__A2 _00747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09460__A1 as2650.stack\[5\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08173__B _02494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10070__A2 _03871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07248_ _01096_ _01662_ _01684_ _01685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__07471__B1 _01903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_10_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08015__A2 _02360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07179_ _01014_ _01596_ _01616_ _01617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_133_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09212__B2 _03107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09763__A2 _00683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08566__A3 _02838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10190_ _00863_ _02722_ _00627_ _04340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_133_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07517__B _01866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09515__A2 _00787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07526__A1 _01932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11322__A2 _01696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_21_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_95_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11713_ _00096_ clknet_leaf_133_wb_clk_i as2650.stack\[14\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10833__A1 _03639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06501__A2 _00937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11644_ _00027_ clknet_leaf_36_wb_clk_i as2650.r123\[0\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_19_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11575_ _04161_ _05616_ _05620_ _05621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09451__A1 _02074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08254__A2 _00850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_155_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06382__I _00653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10526_ _04622_ _04638_ _04639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_13_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11221__C _05278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10457_ _05777_ _00687_ _04571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_124_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08006__A2 _02362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11010__A1 _02746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09754__A2 _00730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10388_ _04404_ _04506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06568__A2 _01011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07765__A1 _02102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08962__B1 _03202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11561__A2 _02732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12127_ net80 net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11986__CLK clknet_leaf_77_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08102__I _02423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11313__A2 _05171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11009_ _02349_ _00599_ _05108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07941__I _02280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10521__B1 _01823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08190__A1 _02505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06550_ _00532_ _00991_ _00993_ _00994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__06557__I _00946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_181_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06481_ as2650.cycle\[8\] _00484_ _00925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09690__A1 _02848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08493__A2 _02741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08220_ _02505_ _02531_ _02532_ _02535_ _00142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_60_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08151_ as2650.stack\[8\]\[13\] _02477_ _02483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08245__A2 _00925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07388__I _01822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07102_ _01520_ _01526_ _01540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_105_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10052__A2 _04120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09993__A2 _03963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08082_ _02419_ _02430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_194_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07033_ _01451_ _01284_ _01472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_134_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_161_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11001__A1 _00451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08548__A3 _01021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09745__A2 net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11001__B2 _00866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06559__A2 _00555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11552__A2 _01498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10542__I _04595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08984_ _03000_ _03222_ _02501_ _03223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_192_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07935_ _02161_ _02231_ _02312_ _02158_ _00080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_4919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07508__A1 _01854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09552__B _02561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07866_ _02214_ _02252_ _02257_ _02261_ _00062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_56_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08181__A1 _02329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07851__I _02033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_186_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09605_ _01005_ _03769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_28_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06817_ _01257_ _01123_ _01259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_95_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11373__I _05455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07797_ _02187_ _02208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_84_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08168__B _02494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09536_ _02563_ _03699_ _03700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06748_ _01060_ _01073_ _01083_ _01191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_58_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10815__A1 _00809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09467_ as2650.stack\[5\]\[7\] _03620_ _03612_ _03635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06679_ _00960_ _01121_ _01122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09681__A1 _01254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06495__A1 _00646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08418_ _02693_ _02701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_185_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10291__A2 _02847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09398_ _03555_ _03575_ _03584_ _03586_ _00269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_156_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08349_ _02133_ _02649_ _02254_ _02650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_36_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06247__A1 _00702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07298__I _01733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10043__A2 _03976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11240__A1 as2650.stack\[6\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09984__A2 _04000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11360_ as2650.r123_2\[3\]\[2\] _05449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07444__B1 _01877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11240__B2 as2650.stack\[4\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_180_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06798__A2 _01239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10311_ _04327_ _04394_ _04443_ _04444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_11291_ _05200_ _01589_ _05382_ _05383_ _03859_ _05384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_106_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10880__C _03641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10242_ _03797_ _04387_ _04389_ _00310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_3_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07747__A1 _02051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11543__A2 _05162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10173_ _04306_ _04322_ _04323_ _04324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__06151__B _00609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_74_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_170_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06722__A2 _00592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06377__I _00755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05930__B1 _05782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10806__A1 _04875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08475__A2 _02747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09672__A1 _03819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05908__S1 _05736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09688__I _03849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06486__A1 _00862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08592__I _02722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_175_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11627_ _02616_ _04443_ _05666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08227__A2 _02538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10034__A2 _04101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11231__A1 _01431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_155_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11558_ _05600_ _05603_ _05604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_171_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07986__A1 net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_176_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07986__B2 _00938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10509_ _04621_ _04622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_11489_ _05546_ _00400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_171_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_174_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10362__I _04482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06410__A1 _00511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05981_ _05813_ _00426_ _00436_ _00439_ _00440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_26_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07720_ _02139_ _02140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11298__A1 _01602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08767__I _03021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07651_ _01028_ _02076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
Xclkbuf_0_wb_clk_i wb_clk_i clknet_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__11193__I _01363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10311__B _04443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06713__A2 _01155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07910__A1 as2650.stack\[10\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06602_ _01035_ _01046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07582_ _00948_ _00929_ _02010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_111_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09321_ _02632_ _03527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06533_ as2650.addr_buff\[5\] _00977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_178_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09663__A1 _02846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08466__A2 _02583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09663__B2 _03819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09598__I _01128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09252_ _03467_ _03469_ _03470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__10273__A2 _04408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11470__A1 _04331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07620__B _02047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06464_ _00577_ _00573_ _00580_ _00581_ _00910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_178_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08203_ _02507_ _02522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11142__B _00914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09183_ _03382_ _03403_ _03404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_147_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10537__I _04648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09415__A1 _02730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06395_ _00838_ _00840_ _00841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_33_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07426__B1 _01859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08134_ _02470_ _02471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11222__A1 _03273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08065_ _02415_ _02406_ _02416_ _02417_ _00105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_clkbuf_leaf_33_wb_clk_i_I clknet_4_7_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_161_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07016_ _01138_ _05793_ _05741_ _01455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_150_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09718__A2 _02808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_161_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_102_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06401__A1 _00843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08967_ _01700_ _03192_ _03205_ _03206_ _03207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_130_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_4716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11289__A1 _05238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07918_ _02128_ _02302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_99_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08898_ _03142_ _01261_ _03125_ _03143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_57_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08154__A1 _02329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07849_ as2650.stack\[13\]\[14\] _02052_ _02248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_44_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07901__A1 _02067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06197__I _00655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10860_ _04326_ _04956_ _04374_ _04965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09519_ _02625_ _03683_ _00293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_31_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10791_ net3 _05721_ _04898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_140_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09654__A1 _00805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_164_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_38_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11461__A1 _02901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_61_wb_clk_i clknet_4_14_0_wb_clk_i clknet_leaf_61_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XPHY_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_40_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_72_wb_clk_i_I clknet_4_11_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_36_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09406__A1 _02177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11412_ as2650.stack\[9\]\[3\] _05478_ _05485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_137_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11343_ as2650.stack\[9\]\[7\] _02142_ _05435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_177_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07756__I _02157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_193_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09709__A2 _03743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11274_ as2650.stack\[1\]\[5\] _01934_ _01936_ as2650.stack\[0\]\[5\] _01937_ as2650.stack\[3\]\[5\]
+ _05368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_101_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_175_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11516__A2 _05243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10182__I _04332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10225_ _00702_ _04374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10724__B1 _01822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09590__B1 _03748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10156_ _00906_ _00986_ _04307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06943__A2 _01382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08587__I _02859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10087_ net40 _04067_ _04165_ _04241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_94_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08145__A1 as2650.stack\[8\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11227__B _00847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08696__A2 _02776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_90_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09645__A1 _03797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08448__A2 _02717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10989_ _04897_ _05080_ _04332_ _05089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_43_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06459__A1 _00645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10785__C _04891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11452__A1 _01223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10255__A2 _04388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06835__I _01034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07120__A2 _01555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06180_ _00638_ _00639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07666__I _02089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06570__I _01013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06631__A1 _01060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11507__A2 _04554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09870_ _02611_ _01457_ _04028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_117_wb_clk_i_I clknet_4_2_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10715__B1 _01789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08821_ _00921_ _03067_ _03068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_154_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10191__A1 _00734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06934__A2 _01109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08752_ _02693_ _03011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05964_ _00422_ _00423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_26_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07703_ _02040_ _02124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_94_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08683_ _01697_ _02955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_113_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_66_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09884__A1 _03975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05895_ _05744_ _05748_ _05749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__08687__A2 _02902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07634_ _02053_ _02060_ _02061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09830__B _03849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10494__A2 _04592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07565_ _01992_ _01993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09636__A1 _03796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08446__B _02718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09304_ _03044_ _03508_ _03512_ _03513_ _00248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__11443__A1 _01295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06516_ as2650.idx_ctrl\[1\] _00960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_22_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11443__B2 as2650.r123\[2\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07496_ _01927_ _01727_ _01928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_146_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08165__C _02494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09235_ _03434_ _03453_ _03454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_167_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06447_ _00576_ _00893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_37_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09166_ _03359_ _03363_ _03386_ _03387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06870__A1 _00439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06378_ _00823_ _00824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_135_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08117_ _02405_ _02454_ _02455_ _02457_ _00117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_09097_ as2650.r0\[1\] _01648_ _03320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08611__A2 _00461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08181__B _02501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07576__I _00925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08048_ _02402_ _02386_ _02403_ _02404_ _00101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__10216__B _03755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05976__A3 _00431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_172_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09791__I net34 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08375__A1 _02198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10010_ _04131_ _03976_ _04165_ _04166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_62_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09999_ _03873_ _04134_ _04155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_114_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_5247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05824__I _05677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08127__A1 _02415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11961_ _00330_ clknet_leaf_15_wb_clk_i as2650.ins_reg\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_57_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09875__A1 _02861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_178_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11131__B1 _05226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_56_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10912_ _04432_ _05002_ _05015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_151_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09740__B _03793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10485__A2 _02039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11892_ _00261_ clknet_leaf_95_wb_clk_i as2650.stack\[3\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10843_ _03665_ _04948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_183_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11434__A1 _05697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07638__B1 _02061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10774_ _02125_ _04880_ _04881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__09031__I _01203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07102__A2 _01526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06861__A1 _01297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06861__B2 _01299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06613__A1 _01007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11326_ net77 _05245_ _05418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_180_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11257_ _00775_ _01501_ _05349_ _05350_ _03813_ _05351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_136_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08366__A1 _02525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10208_ _04352_ _04357_ _04358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_11188_ _03761_ _01303_ _05202_ _05284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_136_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_171_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10139_ _04150_ _04168_ _04291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_95_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08118__A1 _02376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08110__I _02086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_149_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08669__A2 _01141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10476__A2 _04587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10796__B _04897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_189_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10228__A2 _00450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11425__A1 _02184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07350_ _01731_ _01786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06301_ _00572_ _00745_ _00752_ _00010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_176_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07281_ _00838_ _01716_ _01717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_149_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09020_ _03250_ _03251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06232_ _00498_ _00686_ _00689_ _00620_ _00690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_34_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08780__I _02066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06163_ as2650.cycle\[13\] _00622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_172_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06604__A1 _01043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10400__A2 _04480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06094_ _00539_ _00547_ _00552_ _00553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_176_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_171_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09922_ _04078_ _03888_ _03769_ _04079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__06080__A2 _00534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08357__A1 as2650.stack\[3\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09853_ _03975_ _02955_ _04012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10164__A1 _00938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08804_ as2650.stack\[8\]\[7\] _03035_ _03021_ _03052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09784_ _02852_ _03147_ _03851_ _03895_ _03896_ _03944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_06996_ _01435_ _01436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08109__A1 as2650.stack\[0\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08020__I _02128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08735_ _02997_ _02998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05947_ _05797_ _05800_ _05801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_85_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09857__A1 _00629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11113__B1 _05154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08666_ _05695_ _00493_ _02827_ _02938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_96_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10467__A2 _04531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05878_ _05731_ _05732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_187_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07617_ _02044_ _02045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_1728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08597_ _02867_ _02869_ _02870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_26_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11416__A1 _03509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07548_ _01622_ _01911_ _01718_ _01977_ _01978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__05894__A2 _05746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10624__C1 as2650.stack\[10\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07479_ _01717_ _01911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09218_ _03396_ _03436_ _03437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__06843__A1 _01150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10490_ _04584_ _04602_ _04603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_154_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09149_ _03352_ _03370_ _03371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_154_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05819__I _05672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08596__A1 _02346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08596__B2 _01687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_194_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_136_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11111_ _05165_ _05209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_85_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08348__A1 _02648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_5000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11042_ _02819_ _01032_ _05139_ _05140_ _05141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_5011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10155__A1 _03687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11352__B1 _05434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_5044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10170__A4 _04320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_4376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11944_ _00313_ clknet_leaf_63_wb_clk_i as2650.addr_buff\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08865__I _03057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08520__A1 _02780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11875_ _00244_ clknet_leaf_91_wb_clk_i as2650.stack\[2\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_44_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10826_ _04668_ _04931_ _04771_ _04932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11407__A1 _02364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12039__D _00408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10757_ _00521_ _04857_ _04861_ _04864_ _04865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_105_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06834__A1 _01269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_146_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10688_ _04764_ _04766_ _04795_ _04797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_125_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09784__B1 _03851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_154_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10394__A1 _02837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11309_ as2650.stack\[9\]\[6\] _05171_ _05172_ as2650.stack\[11\]\[6\] _05402_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_99_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08339__A1 as2650.stack\[4\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07944__I _02277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10370__I _04482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06850_ _01290_ _01291_ _00967_ _01292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_110_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09551__A3 _03714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06781_ _01107_ _01223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09839__A1 _03995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08520_ _02780_ _02787_ _02792_ _02793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__10449__A2 _00827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08775__I _02466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08451_ _01724_ _02724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_184_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07402_ as2650.stack\[9\]\[9\] _01830_ _01827_ as2650.stack\[8\]\[9\] as2650.stack\[11\]\[9\]
+ _01836_ _01837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_168_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06295__I _00746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08382_ _02672_ _02667_ _02671_ _02674_ _00165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__09067__A2 _03257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11742__CLK clknet_leaf_116_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07333_ _01768_ net73 _01769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_91_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10746__S _04608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08814__A2 _00941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08724__B _02969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06825__A1 _05745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06825__B2 _05739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07264_ _01046_ _01700_ _01040_ _01701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__10621__A2 _01815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09003_ _02989_ _02495_ _03216_ _03237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06215_ _00464_ _00661_ _00671_ _00673_ _00525_ _00674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_07195_ _01541_ _01552_ _01632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_121_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06146_ _00459_ _00605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_30_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10385__A1 _01460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06077_ _00535_ _00536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_99_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_67_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09905_ _04023_ _03959_ _04062_ _04063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__10137__A1 _04102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07002__A1 _01430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_59_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09836_ _03793_ _00723_ _03995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_101_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_47_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08750__A1 _02452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06979_ as2650.holding_reg\[4\] _00830_ _01419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_132_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09767_ _02082_ _03879_ _03927_ _03878_ _03928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_73_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08718_ _02710_ _02985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09698_ _03774_ _03841_ _03858_ _03859_ _03860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_27_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08502__A1 _02749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_2248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08649_ as2650.stack\[15\]\[7\] _01809_ _01814_ as2650.stack\[13\]\[7\] _02921_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_55_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_19_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_11660_ _00043_ clknet_leaf_1_wb_clk_i as2650.stack\[11\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_168_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_165_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07069__A1 _01265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10611_ _03960_ _04721_ _04722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11591_ _05608_ _05606_ _05632_ _05634_ _05635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_195_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08805__A2 _03041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10883__C _04986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10073__B1 _04224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06816__A1 _01255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10542_ _04595_ _04654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_195_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_194_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10473_ _00698_ _04586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_100_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10376__A1 _03148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07241__A1 _01461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08584__A4 _02856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07792__A2 _02197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11025_ _02763_ _02766_ _05116_ _05123_ _05124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__10679__A2 _04701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09533__A3 _03695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08741__A1 _02976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11628__A1 _04444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11765__CLK clknet_leaf_80_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11235__B _05321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11927_ _00296_ clknet_leaf_63_wb_clk_i net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_185_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10851__A2 _04228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11858_ _00227_ clknet_leaf_32_wb_clk_i as2650.r123_2\[0\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_183_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10809_ _04913_ _04914_ _04915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_159_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11789_ _00172_ clknet_4_2_0_wb_clk_i as2650.stack\[1\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_158_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07939__I _02278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06807__A1 _01094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_186_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10603__A2 _04587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10365__I _04480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06000_ as2650.prefixed _00459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_86_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_154_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09221__A2 _02233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06035__A2 _00493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08980__A1 _02143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07951_ as2650.stack\[10\]\[11\] _02319_ _02324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_190_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10119__A1 _04255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10314__B _02609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06902_ _01342_ _01333_ _01343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07882_ _02272_ _02146_ _02147_ _02273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__11129__C _05174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06338__A3 _00787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07535__A2 _01912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09621_ _03732_ _03720_ _03785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06833_ _01274_ _01045_ _01036_ _01275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_110_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11619__A1 _02050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09552_ _02581_ _02584_ _02561_ _03716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06764_ _01106_ _01207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_168_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05922__I _05775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08503_ _02729_ _02736_ _02744_ _02775_ _02776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_102_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09483_ _00973_ _03650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_38_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11095__A2 _00874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06695_ _01120_ _01138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_129_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08434_ as2650.stack\[15\]\[9\] _02712_ _02713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__05849__A2 _05690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08365_ as2650.stack\[3\]\[13\] _02655_ _02661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_20_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08799__A1 as2650.stack\[8\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_1585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07316_ _01751_ _01752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08296_ _02565_ _02587_ _02604_ _02605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_164_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09460__A2 _03615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07247_ _01059_ _01673_ _01681_ _01092_ _01683_ _01684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XANTENNA__07471__A1 _01893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_192_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07178_ _01598_ _01264_ _01014_ _01615_ _01616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_49_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09212__A2 _03342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10358__A1 _03649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07223__A1 _01029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06129_ _00587_ _00588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_106_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07584__I _00928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_86_wb_clk_i clknet_4_2_0_wb_clk_i clknet_leaf_86_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__08971__A1 _01696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10224__B _03649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_15_wb_clk_i clknet_4_5_0_wb_clk_i clknet_leaf_15_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_59_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09515__A3 _03678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11788__CLK clknet_leaf_85_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09819_ _01434_ _03978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output32_I net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_160_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11712_ _00095_ clknet_leaf_1_wb_clk_i as2650.stack\[14\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10833__A2 _01800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11643_ _00026_ clknet_leaf_32_wb_clk_i as2650.r123\[0\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_180_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06663__I _01106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11574_ _00427_ _02813_ _05619_ _03661_ _05620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_126_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09451__A2 _03617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08254__A3 _02550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_168_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_167_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07462__A1 as2650.stack\[2\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10525_ _04630_ _04637_ _04638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_6_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10456_ _04225_ _04570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10349__A1 _00670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11546__B1 _05592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11010__A2 _00502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10387_ net47 _04487_ _04505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_123_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12126_ net80 net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08962__A1 _01563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07765__A2 _02172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11561__A3 _00613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_191_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10134__B _03781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07517__A2 _01944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08714__A1 _02399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11008_ _05102_ _05106_ _05107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_93_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08714__B2 _02982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10521__B2 as2650.stack\[14\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_146_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06774__S net51 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06480_ _05714_ _05728_ _00924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09690__A2 _01286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07669__I net60 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08150_ _02325_ _02480_ _02481_ _02482_ _00125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_187_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10588__A1 _02071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07101_ _01537_ _01525_ _01538_ _01539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07453__A1 _01295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08081_ _02323_ _02420_ _02424_ _02429_ _00109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_174_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_140_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_147_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07032_ _01459_ _01137_ _01470_ _01471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_175_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_3_0_0_wb_clk_i clknet_0_wb_clk_i clknet_3_0_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__07205__A1 _01547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06559__A3 _00973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08953__A1 _01611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11930__CLK clknet_leaf_62_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08983_ _02487_ _03222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06964__B1 _01230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10760__A1 _03642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09833__B _03991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07934_ as2650.stack\[11\]\[13\] _02160_ _02312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_4909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08705__A1 _02384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08705__B2 _02975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07865_ as2650.stack\[12\]\[10\] _02260_ _02261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__10512__A1 _02907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10698__C _02824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09604_ _02844_ _03767_ _03768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_99_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08181__A2 _02500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06816_ _01255_ _01256_ _01257_ _01258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_42_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07796_ _02206_ _02207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_83_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06747_ _00885_ _00515_ _01189_ _01190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_09535_ _00852_ _02588_ _03699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_97_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_133_wb_clk_i clknet_4_1_0_wb_clk_i clknet_leaf_133_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_64_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09466_ _02184_ _03617_ _03634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06678_ _01009_ _01121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__10815__A2 _04152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09681__A2 _01258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_62_wb_clk_i_I clknet_4_14_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06495__A2 _00938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08417_ _02689_ _02700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07692__A1 as2650.stack\[13\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07800__C _02210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09397_ as2650.stack\[6\]\[2\] _03585_ _03582_ _03586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_178_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08348_ _02648_ _02144_ _02649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_177_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10579__A1 _04626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10219__B _04349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06247__A2 _00703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11240__A2 _02387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08279_ _00660_ _00848_ _02574_ _02588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_138_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10310_ _01927_ _04439_ _04443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_193_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11290_ _03761_ _01619_ _05202_ _05383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_125_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10241_ _04186_ _04388_ _04389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05827__I _05680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10172_ _02561_ _02563_ _02594_ _03695_ _04323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_117_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10751__A1 _04023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10503__A1 _02846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08172__A2 _02497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07263__B _01031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06658__I _01101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06183__A1 _00641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10401__C _04506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06722__A3 _01092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05930__A1 _05781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_186_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_147_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08873__I _03057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10806__A2 _04789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xwrapped_as2650_160 la_data_out[49] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_187_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08475__A3 _00598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06486__A2 _00929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11513__B _05192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11626_ _05674_ _04394_ _02340_ _05665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_168_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11231__A2 _05138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11557_ _00754_ _04621_ _05601_ _02740_ _05602_ _05603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_156_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07986__A2 _02340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10508_ _00929_ _02727_ _04621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11488_ as2650.r123\[3\]\[1\] _05546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11953__CLK clknet_leaf_20_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_195_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10990__A1 _04863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10439_ _04545_ _04552_ _04553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_154_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_107_wb_clk_i_I clknet_4_3_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08113__I _02423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06410__A2 _00765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05980_ _00437_ _00438_ _00439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11298__A2 _02960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09360__A1 _02074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07650_ _02067_ _01998_ _02068_ _02075_ _00032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_65_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06601_ _01044_ _01045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_78_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07910__A2 _02293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07581_ _00518_ _02006_ _02007_ _02008_ _02009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_53_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_165_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09112__A1 _03305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09320_ _03520_ _03526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_81_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06532_ as2650.addr_buff\[6\] _00976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_39_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09663__A2 _00683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09251_ _03466_ _03468_ _03469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06463_ _00509_ _00586_ _00901_ _00908_ _00909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_142_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11470__A2 _00950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08202_ _02226_ _02521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09182_ _03385_ _03402_ _03403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_193_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06394_ _00503_ _00839_ _00667_ _00840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_105_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09415__A2 _02580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08133_ _01991_ _02144_ _02470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_146_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07426__B2 as2650.stack\[5\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08064_ _02302_ _02258_ _02385_ _02417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_50_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_11_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10981__A1 _04595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09179__A1 _03395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07015_ _05802_ _05807_ _05810_ _01454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_134_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09718__A3 _03879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08926__A1 _01431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10733__A1 as2650.ivec\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_192_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_142_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10733__B2 _04793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08966_ _02932_ _03114_ _03192_ _03206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_4706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11289__A2 _04081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07917_ as2650.stack\[10\]\[7\] _02293_ _02301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_4739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08897_ _03122_ _03132_ _03140_ _03141_ _03142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_116_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08154__A2 _02480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08179__B _02501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09351__A1 _03542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_186_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06165__A1 _00553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07848_ _02053_ _02231_ _02247_ _02047_ _00058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_17_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07779_ _02190_ _02191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__11826__CLK clknet_leaf_106_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09518_ _03671_ _03672_ _03682_ _03683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_140_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08693__I _02964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10790_ _03746_ _04897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09654__A2 _00816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08626__C _01416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_160_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__11461__A2 _02844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09449_ _03550_ _03613_ _03619_ _03622_ _00284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_185_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_16_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09406__A2 _03579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11976__CLK clknet_leaf_75_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11411_ _03555_ _05473_ _05483_ _05484_ _00384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_123_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09738__B _00641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11342_ _05430_ _05433_ _05152_ _05434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_137_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_30_wb_clk_i clknet_4_7_0_wb_clk_i clknet_leaf_30_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__10972__A1 _00522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11273_ as2650.stack\[2\]\[5\] _05225_ _05367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_141_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08917__A1 _01350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10224_ _03686_ _04309_ _03649_ _04373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_171_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10724__A1 as2650.stack\[15\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10724__B2 as2650.stack\[14\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09590__A1 _03737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10155_ _03687_ _03690_ _04306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08868__I _03081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10086_ _02212_ _03788_ _04239_ _04163_ _04240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_59_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08089__B _02431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08145__A2 _02477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09342__A1 _03050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06388__I _00658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09893__A2 _02933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09645__A2 _03803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10988_ _04439_ _05082_ _05087_ _04904_ _05088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__06459__A2 _00904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11452__A2 _03473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_128_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_182_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_188_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07012__I _05802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11609_ _01290_ _05648_ _05651_ _05647_ _05652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_129_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08552__B _02822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07947__I _02213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_195_1927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06851__I _01292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08081__A1 _02323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10373__I _04480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08908__A1 _00439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10715__A1 as2650.stack\[6\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10715__B2 as2650.stack\[5\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08820_ _03060_ _03063_ _03065_ _03066_ _03067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_119_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06395__A1 _00838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10191__A2 _00450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07682__I net61 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05963_ _00420_ _00421_ _00422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_39_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08751_ _02402_ _02996_ _03009_ _03010_ _00198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_57_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10322__B _02353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11849__CLK clknet_4_12_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09333__A1 _03040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07702_ as2650.stack\[13\]\[7\] _02062_ _02123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_187_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05894_ _05745_ _05746_ _05747_ _05739_ _05748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_08682_ _02597_ _02950_ _02953_ _02954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XANTENNA__11140__A1 _04275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08931__I1 _01422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07633_ _02059_ _02060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_26_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08727__B _02969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10976__C _05076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07564_ net73 _01992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_41_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11999__CLK clknet_4_15_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09636__A2 _01118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09402__I _02511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06515_ _00772_ _00958_ _00959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09303_ as2650.stack\[2\]\[5\] _03504_ _03493_ _03513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_110_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07647__A1 _02071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11443__A2 _05502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07495_ _01430_ _01927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_161_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09234_ _03435_ _03452_ _03453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_142_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06446_ _00891_ _00567_ _00892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09165_ _03364_ _03368_ _03386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__06870__A2 _00932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06377_ _00755_ _00823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_194_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_163_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08116_ _02456_ _02425_ _02446_ _02457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_147_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09096_ _01645_ _03317_ _03318_ _03319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_134_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08047_ _02170_ _02392_ _02397_ _02404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_134_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10706__A1 _04397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09572__A1 _00795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08375__A2 _02649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08688__I _02592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06386__A1 _00826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09998_ _04131_ _03867_ _04154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_88_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_5259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08949_ _03176_ _03190_ _00216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_4525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08127__A2 _02454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09324__A1 as2650.stack\[4\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11960_ _00329_ clknet_4_7_0_wb_clk_i as2650.ins_reg\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11047__C _00823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06138__A1 _00594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11131__A1 as2650.stack\[13\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09875__A2 _03850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11131__B2 as2650.stack\[12\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06001__I _05771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10911_ _05006_ _05011_ _05013_ _05014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_3868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07886__A1 _02186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10485__A3 _00804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11891_ _00260_ clknet_leaf_94_wb_clk_i as2650.stack\[3\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_2_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10842_ _04946_ _04947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_96_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__12004__CLK clknet_leaf_120_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05840__I _05693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07638__A1 _02051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10773_ _02115_ _04801_ _04880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_73_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06310__A1 _00757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06861__A2 _01010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11198__A1 _00439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07767__I _02118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08063__A1 as2650.stack\[12\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10945__A1 _04897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10193__I _04341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11325_ _05249_ _03465_ _05417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07810__A1 _01363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07810__B2 _02218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11256_ _04409_ _01458_ _00914_ _05350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_134_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09563__A1 _00804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10207_ _03700_ _03716_ _04354_ _04356_ _04357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_11187_ _05238_ _03147_ _05283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_95_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10173__A2 _04322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10138_ _02225_ _04101_ _04289_ _04290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_67_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09315__A1 as2650.stack\[4\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10069_ _04222_ _04223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_23_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_169_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07877__A1 _02198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10796__C _04902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06846__I _01250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11425__A2 _05480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06300_ _00707_ _00751_ _00752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07280_ _01605_ _01714_ _01715_ _01716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_31_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06301__A1 _00572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06231_ _00688_ _00689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_125_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06852__A2 _01261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07677__I net52 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06162_ _00620_ _00621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_144_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06093_ _00551_ _00552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09921_ _04077_ _04078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06080__A3 _00538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08357__A2 _02655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09554__A1 _03684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09852_ _03975_ _03742_ _03997_ _04009_ _04010_ _04011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_113_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06368__A1 _00739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10164__A2 _02333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08803_ _02381_ _02475_ _03051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08301__I net75 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09783_ _02853_ _03147_ _03943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_112_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06995_ _01434_ _01435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_132_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08109__A2 _02440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09306__A1 _03239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08734_ _02003_ _02437_ _02147_ _02997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_67_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_73_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12027__CLK clknet_leaf_39_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05946_ _05798_ _05786_ _05799_ _05800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_96_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11113__A1 as2650.stack\[4\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11113__B2 as2650.stack\[7\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07868__A1 _02220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05877_ as2650.r0\[5\] _05731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08665_ _02342_ _02335_ _02827_ _02937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_167_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07616_ _02039_ _02041_ _02043_ _02044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__06756__I _01198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08596_ _02346_ _00769_ _02821_ _02868_ _01687_ _02869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_109_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07547_ _01890_ _01974_ _01976_ _01802_ _01977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__11416__A2 _05480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10624__B1 _01818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07478_ _01719_ _01910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08293__A1 _00735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10624__C2 _01876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_194_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08293__B2 _02593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09217_ _05733_ _03393_ _03436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_10_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11611__B _05647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06843__A2 _01284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06429_ _00471_ _00870_ _00874_ _00875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_10_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09148_ _03355_ _03369_ _03370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_120_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08596__A2 _00769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09079_ _01631_ _01655_ _03302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_120_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11110_ _05199_ _05207_ _00824_ _05208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_162_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_172_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11041_ _02812_ _05140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09545__A1 _02556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06359__A1 _00550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07536__B _01735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output62_I net62 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11352__A1 _05413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_5045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_162_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_162_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11943_ _00312_ clknet_leaf_56_wb_clk_i as2650.addr_buff\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_4399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_185_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06666__I _01109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06531__A1 _00542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11874_ _00243_ clknet_leaf_90_wb_clk_i as2650.stack\[2\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_45_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_189_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09042__I _03258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10825_ _04116_ _04930_ _04931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_2997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11407__A2 _05480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_186_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08881__I _03065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08284__A1 _00506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10756_ _04862_ _04863_ _04864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_92_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10091__A1 _04242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_185_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10687_ _04764_ _04766_ _04795_ _04796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_145_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05893__I0 as2650.r123\[1\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08036__A1 _02060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11240__C _05298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10918__A1 _04584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09784__A1 _02852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09926__B _04082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11591__A1 _05608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11308_ _05397_ _05400_ _05265_ _05401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_141_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09645__C _00534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08339__A2 _02636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09536__A1 _02563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11239_ as2650.stack\[5\]\[4\] _05302_ _05163_ as2650.stack\[7\]\[4\] _05334_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_155_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11343__A1 as2650.stack\[9\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07011__A2 _01450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_27_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06780_ _01202_ _01221_ _01222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_97_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09839__A2 _03997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08277__B _02585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06576__I _05776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08450_ _02722_ _02723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_23_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07401_ _01835_ _01836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_51_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08381_ as2650.stack\[2\]\[9\] _02673_ _02674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_91_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_162_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07332_ net70 _01768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08275__A1 _00860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07263_ _01028_ _00427_ _01031_ _01700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__06825__A2 _05767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05884__I0 as2650.r123\[1\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06214_ _00672_ _00673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09002_ as2650.stack\[7\]\[5\] _03220_ _03236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_121_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07194_ _01553_ _01629_ _01630_ _01631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10909__A1 _04391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_191_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06145_ _00600_ _00603_ _00509_ _00604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_195_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06589__A1 _01027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11582__A1 _05138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_172_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07250__A2 _01454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06076_ net6 _00535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09904_ _02745_ _04062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_113_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10137__A2 _04278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07538__B1 _01941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07538__C2 _01870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09835_ _00718_ _03993_ _03994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_115_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11593__S _01685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08750__A2 _03001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09766_ _03917_ _03923_ _03926_ _03927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_58_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06978_ _01094_ _01415_ _01417_ _01418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__07870__I _02256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08717_ _02402_ _02970_ _02983_ _02984_ _00190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_2205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05929_ as2650.r123\[1\]\[1\] as2650.r123\[0\]\[1\] as2650.r123_2\[1\]\[1\] as2650.r123_2\[0\]\[1\]
+ _05705_ _05753_ _05783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
X_09697_ _02889_ _03859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08648_ as2650.stack\[14\]\[7\] _01875_ _01817_ as2650.stack\[12\]\[7\] _02920_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_148_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08579_ net11 _02852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_25_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_74_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__10448__I0 _02038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09797__I net60 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10610_ _04669_ _04673_ _04719_ _04721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XPHY_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_167_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08266__A1 _00886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11590_ _00662_ _05633_ _05634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10073__A1 _04223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_167_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06816__A2 _01256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10073__B2 _04226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10541_ _02069_ _04597_ _04653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_167_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08018__A1 _02181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10472_ _04186_ _03873_ _04585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_10_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09766__A1 _03917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11573__A1 _02834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_123_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07266__B _01132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10471__I _00783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11325__A1 _05249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_150_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_49_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11024_ _02734_ _05118_ _05122_ _05123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_133_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09533__A4 _03696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08741__A2 _02700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08876__I _03062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06752__A1 _01166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11516__B _02570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_4_2_0_wb_clk_i clknet_3_1_0_wb_clk_i clknet_4_2_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_3462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11926_ _00295_ clknet_leaf_62_wb_clk_i net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06396__I _00841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_60_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10300__A2 _04434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11857_ _00004_ clknet_4_12_0_wb_clk_i as2650.cycle\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10808_ _04875_ _04876_ _04914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_158_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11788_ _00171_ clknet_leaf_85_wb_clk_i as2650.stack\[1\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_13_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06807__A2 _01230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10739_ _04229_ _05746_ _04847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_35_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07020__I _05733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10367__A2 _04486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11564__A1 _02076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_192_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09509__A1 _00572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07950_ _02219_ _02323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_9_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10119__A2 _04118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06901_ _01331_ _01342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_122_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07881_ _02271_ _02272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09620_ _03723_ _03725_ _03758_ _03783_ _03784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_110_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06832_ _01273_ _01274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__11331__A4 _05422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07690__I _05682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09551_ _03711_ _03712_ _03714_ _03715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_06763_ _01202_ _01205_ _01206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_55_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10330__B _04343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08502_ _02749_ _02767_ _02774_ _02775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_97_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06694_ _00943_ _01137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_129_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09482_ _03648_ _03649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_110_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08496__A1 _02730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05929__S0 _05705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_52_wb_clk_i_I clknet_4_13_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08433_ _02705_ _02712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05849__A3 _05695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08248__A1 _00470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08364_ _02521_ _02658_ _02659_ _02660_ _00161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_51_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08799__A2 _03026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07315_ _01750_ _01751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11252__B1 _05337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10556__I _04570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08295_ _02588_ _02590_ _02591_ _02603_ _02604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_176_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_192_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07246_ _01341_ _01674_ _01682_ _01498_ _01165_ _01683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_192_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09748__A1 _03876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07177_ _01264_ _01614_ _01615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_121_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10358__A2 _04476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11555__A1 _00773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06128_ _00463_ _05679_ _00587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08420__A1 _02680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_1384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06059_ _00513_ _00517_ _00518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_156_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11307__A1 _05364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09515__A4 _03679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09818_ _00748_ _03977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_100_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_91_wb_clk_i_I clknet_4_8_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06734__A1 _00885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_55_wb_clk_i clknet_4_12_0_wb_clk_i clknet_leaf_55_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_143_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09749_ _03861_ _03840_ _03909_ _03910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_41_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_95_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08487__A1 _02759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output25_I net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07105__I _01542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11711_ _00094_ clknet_leaf_133_wb_clk_i as2650.stack\[14\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08645__B _01844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11642_ _00025_ clknet_leaf_37_wb_clk_i as2650.r123\[0\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08239__A1 _00524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09320__I _03520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11243__B1 _05172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11573_ _02834_ _02819_ _05618_ _05140_ _05619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__06165__B _00623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10524_ _01845_ _04633_ _04636_ _04637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_168_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07462__A2 _01865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10455_ _04428_ _04564_ _04567_ _04568_ _04569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__09476__B _03642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_182_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10349__A2 _03673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11546__B2 _02621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08411__A1 _02672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10386_ _03279_ _04483_ _04503_ _04504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11010__A3 _03638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06612__C _01055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12125_ net80 net17 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08962__A2 _03177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11561__A4 _05131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_156_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06973__A1 _01392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11732__CLK clknet_leaf_108_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08714__A2 _02970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11007_ _02568_ _02731_ _02739_ _05105_ _05106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_78_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06725__A1 _00434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10521__A2 _01810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_93_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10150__B _04301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08478__A1 _02577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_185_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10285__A1 _04419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11909_ _00278_ clknet_leaf_75_wb_clk_i as2650.ivec\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07150__A1 _01327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08555__B _02723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09690__A3 _03851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09978__A1 _04131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_186_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_147_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10588__A2 _04531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07100_ _01393_ _01201_ _01523_ _01538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_147_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08080_ as2650.stack\[0\]\[11\] _02427_ _02429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_147_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08650__A1 _01764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07031_ _01460_ _01140_ _01469_ _00944_ _01470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_122_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11537__A1 _05579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06559__A4 _01002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08982_ as2650.stack\[7\]\[0\] _03220_ _03221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_157_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06964__B2 _01235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10760__A2 _04859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07933_ _02161_ _02227_ _02311_ _02158_ _00079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_111_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09902__A1 _00896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08705__A2 _02970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07864_ _02250_ _02260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_29_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09603_ _03766_ _03092_ _03767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06815_ _01008_ _01009_ _01257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_110_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07795_ _01204_ _02191_ _02192_ _02205_ _02206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_37_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09534_ _03687_ _03690_ _03693_ _03697_ _03698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_06746_ _01184_ _01187_ _01186_ _01189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_37_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08469__A1 _00883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10995__B _05093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10276__A1 _04400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09465_ _03568_ _03627_ _03632_ _03633_ _00289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06677_ _00429_ _01120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_145_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07141__A1 _01059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09681__A3 _01260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08416_ _02678_ _02690_ _02694_ _02699_ _00174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_51_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06764__I _01106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_145_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07692__A2 _02062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09396_ _03576_ _03585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10028__A1 _04181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10286__I _04422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08347_ _02135_ _02648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_177_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_22_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_102_wb_clk_i clknet_4_9_0_wb_clk_i clknet_leaf_102_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__07444__A2 _01874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08278_ _02566_ _02569_ _02579_ _02586_ _02587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_138_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07229_ _01029_ _00991_ _01665_ _01486_ _01666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_101_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11528__A1 _04462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07595__I _02022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10240_ _04385_ _04388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11755__CLK clknet_leaf_81_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10200__A1 _00548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10171_ _00723_ _04308_ _04310_ _04312_ _04321_ _04322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_105_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06955__A1 _05806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10751__A2 _03733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06004__I as2650.ins_reg\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11992__D _00361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06939__I _01378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_170_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10503__A2 _04586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11161__C1 as2650.stack\[6\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05915__C1 _05768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10267__A1 _03673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11464__B1 _05521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xwrapped_as2650_150 io_oeb[36] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_128_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07132__A1 _05748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_161 la_data_out[51] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_42_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08475__A4 _00603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11513__C _02608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11625_ _05662_ _05664_ _00418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_15_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11216__B1 _05178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08632__A1 _00958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11556_ _00736_ _02841_ _00950_ _02735_ _05602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_156_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10507_ _04534_ _04620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_11487_ _05545_ _00399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_183_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11519__A1 _02777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10438_ _01775_ _04548_ _04551_ _04552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__07199__A1 _05765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10369_ _04482_ _04490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_151_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09426__S _03604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06410__A3 _00855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12039_ _00408_ clknet_leaf_19_wb_clk_i as2650.ins_reg\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06849__I _00957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_66_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06600_ _00923_ _00946_ _00927_ _00931_ _01044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_25_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07580_ _01603_ _02008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_19_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06531_ _00542_ _00974_ _00975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_94_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07123__A1 _01539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_0_wb_clk_i clknet_4_1_0_wb_clk_i clknet_leaf_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_80_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09250_ _01663_ _02234_ _03468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_90_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06584__I net50 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06462_ _00902_ _00907_ _05677_ _00749_ _00908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_107_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08871__A1 _01146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07674__A2 _02097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08201_ _02519_ _02508_ _02512_ _02520_ _00138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__06882__B1 _01322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09181_ _03387_ _03401_ _03402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_06393_ _00590_ _05695_ _00839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_187_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08132_ as2650.stack\[8\]\[8\] _02467_ _02469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_119_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07426__A2 _01858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08623__A1 _02776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10430__A1 _04540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08063_ as2650.stack\[12\]\[7\] _02396_ _02416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_146_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09179__A2 _03399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07014_ _01451_ _01452_ _01453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__08304__I _02612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06937__A1 _05752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10733__A2 _04470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08965_ _05796_ _03151_ _03205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_4707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_170_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07916_ _02113_ _02292_ _02299_ _02300_ _00073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_4729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08896_ _01286_ _03063_ _03141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_130_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_57_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07847_ as2650.stack\[13\]\[13\] _02052_ _02247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_17_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07778_ _02020_ _02190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_140_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09517_ _02726_ _03673_ _03677_ _03681_ _03682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_06729_ _01065_ _00989_ _01135_ _01172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_25_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07114__A1 _01547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_77_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09448_ as2650.stack\[5\]\[1\] _03620_ _03621_ _03622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08862__A1 _01102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_181_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09379_ _02121_ _03571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_8_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11410_ _02074_ _05480_ _05481_ _05484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_149_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08614__A1 _01422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11341_ _05216_ _05431_ _05432_ _05433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_193_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_180_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07539__B _01735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06443__B _00877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10972__A2 _05059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08214__I _02529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11272_ as2650.stack\[5\]\[5\] _05302_ _05303_ as2650.stack\[7\]\[5\] as2650.stack\[6\]\[5\]
+ _05296_ _05366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_152_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_181_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10223_ _00565_ _00700_ _00741_ _04348_ _04372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_152_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_180_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_165_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10724__A2 _04822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_70_wb_clk_i clknet_4_11_0_wb_clk_i clknet_leaf_70_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_133_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09590__A2 _03738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10154_ _03699_ _04304_ _04305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_121_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10085_ _04212_ _04221_ _04238_ _04161_ _04239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_121_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11524__I1 _02001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09045__I _01905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10488__A1 _04596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09342__A2 _03533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_188_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08884__I _03104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10987_ _04400_ _05083_ _05086_ _00586_ _02901_ _05087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_62_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_128_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08853__A1 _00606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11608_ _02778_ _04786_ _05650_ _05651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_160_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08552__C _02824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11539_ _05576_ _05586_ _04501_ _05587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_128_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08081__A2 _02420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06092__A1 _00549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08908__A2 _03058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_171_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10715__A2 _04542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07963__I _02331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06395__A2 _00840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07592__A1 _00861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08750_ _02452_ _03001_ _03005_ _03010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_85_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05962_ _05719_ _05754_ _05755_ _05707_ _00421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_117_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10479__A1 _00809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07701_ _02121_ _02122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09333__A2 _03533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08681_ _02951_ _02952_ _02335_ _02827_ _02953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_66_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05893_ as2650.r123\[1\]\[6\] as2650.r123\[0\]\[6\] as2650.r123_2\[1\]\[6\] as2650.r123_2\[0\]\[6\]
+ _05684_ _05713_ _05747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_65_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11140__A2 _01261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07632_ _02057_ _02041_ _02058_ _02059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_93_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07912__B _02269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08794__I _02101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09097__A1 as2650.r0\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07563_ _01990_ _01991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09636__A3 _01158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09302_ _02376_ _03502_ _03512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_55_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06514_ _00663_ _00461_ _00958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08844__A1 _01019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07494_ _01916_ _01919_ _01925_ _01799_ _01926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_126_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09233_ _03447_ _03451_ _03452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__10651__A1 _05673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06445_ _00557_ _00545_ _00891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09839__B _03776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10992__C _04364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_4_15_0_wb_clk_i clknet_3_7_0_wb_clk_i clknet_4_15_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_21_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09164_ _03383_ _03384_ _03385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_148_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06376_ _00731_ _00822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_120_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08115_ _02096_ _02456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10403__A1 _02602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09095_ _01546_ _01651_ _03318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08046_ as2650.stack\[12\]\[3\] _02390_ _02403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_135_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_176_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_118_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09572__A2 _03731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08375__A3 _02254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09997_ _03734_ _04152_ _04153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07806__C _02210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07583__A1 _00878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06386__A2 _00827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08948_ _01530_ _03177_ _03189_ _03099_ _03190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_4504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06489__I _00932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09324__A2 _03521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08879_ _03070_ _03125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_91_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11131__A2 _02142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10910_ _04609_ _05012_ _04724_ _05013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_29_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06689__A3 _01131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11890_ _00259_ clknet_leaf_95_wb_clk_i as2650.stack\[3\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_56_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11943__CLK clknet_leaf_56_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10841_ _04167_ _04945_ _04946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_71_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10890__A1 _04948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10772_ _00782_ _04879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07638__A2 _01998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06310__A2 _00696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08653__B _02776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10474__I _04586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10945__A2 _05046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11324_ _00775_ _01685_ _05414_ _05415_ _03813_ _05416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_114_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11255_ _04129_ _01474_ _05349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09012__A1 _05696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08879__I _03070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10206_ _03692_ _02594_ _03676_ _04355_ _04356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XANTENNA__09563__A2 _02865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11186_ _00680_ _05282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_121_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10137_ _04102_ _04278_ _04288_ _04289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_121_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06399__I _00844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09315__A2 _03521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10068_ net66 _04222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_82_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08523__B1 _02795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_91_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07877__A2 _02136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_47_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10881__A1 _04794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09079__A1 _01631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_149_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07023__I _01461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_182_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_188_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06301__A2 _00745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06230_ _00687_ _00688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_164_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06862__I _01302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11189__A2 _01350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06161_ _00529_ _00584_ _00619_ _00620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_69_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_1714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_195_1725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06065__A1 _00487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10936__A2 _05033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06092_ _00549_ _00550_ _00551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_102_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09920_ _04076_ _04077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11816__CLK clknet_leaf_111_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09003__A1 _02989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08789__I _02090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06811__B _01227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07693__I net62 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_193_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09851_ _03870_ _02612_ _03743_ _04010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_119_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10333__B _04343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06368__A2 _00625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10164__A3 _04314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08802_ _02121_ _03050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_140_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09782_ _02859_ _03803_ _00534_ _03942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_140_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06994_ net12 _01434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08733_ _02995_ _02996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09306__A2 _02673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05945_ _05735_ _05740_ _05799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_100_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_54_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11113__A2 _05210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10987__C _02901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08664_ _02928_ _02929_ _02935_ _02936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_94_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05876_ _05716_ _05722_ _05729_ _05730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_27_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07868__A2 _02252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07615_ _01100_ _02042_ _02043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__10872__A1 _04199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08595_ _02834_ _00769_ _02868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_42_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06540__A2 _00981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07546_ _01975_ _01727_ _01976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08817__A1 _02089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10624__A1 as2650.stack\[9\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10624__B2 as2650.stack\[8\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07477_ as2650.r123\[0\]\[4\] _01909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__08293__A2 _00490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09216_ _03426_ _03428_ _03435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06428_ _00873_ _00874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09147_ _03364_ _03368_ _03369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_135_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06359_ _00550_ _00692_ _00807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10927__A2 _04293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09078_ _01634_ _01654_ _03301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_159_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08596__A3 _02821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08029_ _01999_ _02001_ _02388_ _02023_ _02389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_151_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08699__I _02969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11040_ _05129_ _01111_ _05137_ _05138_ _05139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_5002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06359__A2 _00692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_104_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11352__A2 _05427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_77_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output55_I net90 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11942_ _00311_ clknet_leaf_56_wb_clk_i as2650.addr_buff\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_4378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05851__I as2650.ins_reg\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10469__I _04581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11873_ _00242_ clknet_leaf_40_wb_clk_i as2650.r123_2\[2\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06531__A2 _00974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10824_ _04929_ _04899_ _00698_ _04930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_2987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10615__A1 _04720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10755_ _04400_ _00699_ _04105_ _04863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09481__A1 _02806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08284__A2 _02004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07778__I _02020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_186_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10686_ _01464_ _05737_ _04795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_173_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05893__I1 as2650.r123\[0\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08036__A2 _02263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11040__A1 _05129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09784__A2 _03147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07795__A1 _01204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11307_ _05364_ _05398_ _05399_ _05400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__07795__B2 _02205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11989__CLK clknet_leaf_75_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08402__I _02688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11238_ _05331_ _05332_ _05333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09536__A2 _03699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11343__A2 _02142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11169_ _01782_ _05266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_23_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07462__B _01866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08898__I1 _01261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10854__A1 _04590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07180__C1 _01593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07400_ _01809_ _01835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08380_ _02665_ _02673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10606__A1 _05673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07331_ as2650.stack\[2\]\[8\] _01747_ _01766_ _01767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_36_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08275__A2 _02583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06592__I _01035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07262_ _01697_ _00934_ _01145_ _01698_ _01699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_104_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07483__B1 _01856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_176_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_192_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09001_ _03040_ _03233_ _03234_ _03235_ _00223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06213_ _00608_ _00672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__05884__I1 as2650.r123\[0\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07193_ _01555_ _01557_ _01630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10909__A2 _03873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06038__A1 _05676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06144_ _00494_ _00602_ _00603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_121_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06589__A2 _01032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11582__A2 _04446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10842__I _04946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06075_ _00533_ _00534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07637__B _02063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05936__I _05779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_99_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09903_ _04058_ _04060_ _03968_ _04061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09527__A2 _00579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08312__I _02571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09834_ _03983_ _03984_ _03990_ _03992_ _03993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xclkbuf_leaf_127_wb_clk_i clknet_4_1_0_wb_clk_i clknet_leaf_127_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_101_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_81_wb_clk_i_I clknet_4_8_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06210__A1 _05704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09765_ _00689_ _03903_ _03924_ _03925_ _03926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_101_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06977_ _00885_ _00766_ _01416_ _01417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_189_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11098__A1 _05129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08716_ _02452_ _02974_ _02979_ _02984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05928_ as2650.r123\[2\]\[1\] as2650.r123_2\[2\]\[1\] _05753_ _05782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_09696_ _03793_ _03855_ _03857_ _03771_ _00551_ _03858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_6_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10289__I _04422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10845__A1 _02195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08647_ as2650.stack\[10\]\[7\] _02909_ _01764_ _02919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_2239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08502__A3 _02774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05859_ _05712_ _05713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07710__A1 _02122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08578_ _02850_ _02851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_14_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_39_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_23_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07529_ _01874_ _01959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07069__A3 _01361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08266__A2 _00686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09463__A1 as2650.stack\[5\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10073__A2 _03752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10540_ _04651_ _04652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_195_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10471_ _00783_ _04584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08018__A2 _02202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06029__A1 _00487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11022__A1 _00864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11995__D _00364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11573__A2 _02819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11325__A2 _03465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11023_ _05120_ _05121_ _02742_ _05122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_77_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06201__A1 _00648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_65_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11089__A1 _01102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10199__I _02572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10836__A1 as2650.ivec\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11925_ _00294_ clknet_leaf_62_wb_clk_i net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10836__B2 _04934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11856_ _00003_ clknet_leaf_66_wb_clk_i as2650.cycle\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10807_ _02194_ _04913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_32_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11787_ _00170_ clknet_leaf_85_wb_clk_i as2650.stack\[2\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_126_wb_clk_i_I clknet_4_0_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09454__A1 _02087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06268__A1 _00549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11261__A1 _02724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10738_ _04844_ _04846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_185_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07301__I _01736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10669_ _04777_ _04778_ _01775_ _04779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_127_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_173_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12017__CLK clknet_leaf_101_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11013__A1 _00722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07768__A1 _02181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_9_wb_clk_i_I clknet_4_4_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10119__A3 _04120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11316__A2 _05408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06900_ _01086_ _01341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07880_ _01762_ _02271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_60_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08193__A1 as2650.stack\[6\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06831_ _01272_ _01273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_95_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06743__A2 _01068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09550_ _02552_ _03713_ _00607_ _00956_ _03714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_06762_ _01203_ _01112_ _01204_ _01101_ _01205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_110_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10330__C _04458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08501_ _00853_ _02768_ _02771_ _02773_ _02774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__10827__A1 _04668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09481_ _02806_ _03647_ _03648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_149_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09693__A1 _03848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06693_ _01135_ _01136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08496__A2 _02341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05929__S1 _05753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08432_ _02663_ _02707_ _02708_ _02711_ _00178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_63_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08363_ as2650.stack\[3\]\[12\] _02655_ _02660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_71_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09445__A1 _02284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06259__A1 _00714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07314_ _01749_ _01750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_162_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11252__A1 _00757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08294_ _02594_ _02601_ _02602_ _02603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_164_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07245_ _01675_ _01682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_118_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_176_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05867__S _05713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11004__A1 _03243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_191_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09748__A2 net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_180_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07176_ _01599_ _01307_ _01613_ _01614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07759__A1 _02174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11555__A2 _01090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06127_ _00585_ _00586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_160_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08420__A2 _02700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10505__C _04333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06431__A1 _00617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06058_ _00449_ _00516_ _00517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_8_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10515__B1 _02909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08977__I _02492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07881__I _02271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09817_ _03719_ _03976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11617__B _04430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06497__I _00478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09748_ _03876_ net10 _03909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_132_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10818__A1 _04709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09679_ _03838_ _03840_ _03841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_54_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09684__A1 _03842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08487__A2 _01711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11710_ _00093_ clknet_leaf_133_wb_clk_i as2650.stack\[14\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_42_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_95_wb_clk_i clknet_4_9_0_wb_clk_i clknet_leaf_95_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_54_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10294__A2 _04429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output18_I net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_187_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11641_ _00024_ clknet_leaf_36_wb_clk_i as2650.r123\[0\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08239__A2 _00758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09436__A1 _01980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_145_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11243__A1 as2650.stack\[13\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11572_ _05138_ _04417_ _05617_ _05618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__11243__B2 as2650.stack\[15\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10523_ _01765_ _04634_ _04635_ _04636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_183_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09739__A2 _03898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10454_ _04156_ _00520_ _00894_ _04568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_87_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11546__A2 _05565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10349__A3 _02741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10482__I _00443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10385_ _01460_ _04484_ _04503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08411__A2 _02690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11010__A4 _05108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12124_ net80 net16 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06422__A1 _00865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_61_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11006_ _00766_ _00648_ _00870_ _05104_ _05105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_77_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10809__A1 _04913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_52_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11908_ _00277_ clknet_leaf_71_wb_clk_i as2650.ivec\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11482__A1 _04652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_163_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11839_ _00222_ clknet_leaf_97_wb_clk_i as2650.stack\[7\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11234__A1 _03815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07030_ _01462_ _01046_ _01039_ _01468_ _01469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_173_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_162_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06661__A1 _01103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_161_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_177_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06413__A1 _00831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08981_ _03219_ _03220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_9_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_170_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07932_ as2650.stack\[11\]\[12\] _02307_ _02311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_151_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07915__B _02269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09902__A2 _04043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07863_ _02207_ _02252_ _02257_ _02259_ _00061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_96_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06716__A2 _01158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10341__B _04466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07913__A1 _02102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11170__B1 _02002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06814_ _01138_ _00432_ _01227_ _01256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_09602_ _00991_ _03766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07794_ _02204_ _02205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_37_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09533_ _02585_ _02578_ _03695_ _03696_ _03697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_168_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06745_ _01184_ _01186_ _01187_ _01188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_1920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08469__A2 _00832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09666__B2 _03827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10276__A2 _00822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09464_ _02119_ _02536_ _03612_ _03633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06676_ _01118_ _01119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_36_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08415_ as2650.stack\[1\]\[11\] _02697_ _02699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_58_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09395_ _02167_ _02522_ _03584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11225__A1 _03948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08346_ as2650.stack\[3\]\[8\] _02645_ _02647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_149_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09969__A2 _01695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08037__I _02389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_20_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08277_ _02581_ _02584_ _02585_ _02586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_20_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07228_ _01664_ _00990_ _01665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11528__A2 _05575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07159_ _01569_ _01597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06404__A1 _00514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10170_ _03677_ _04316_ _04318_ _04320_ _04321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_154_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_154_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08157__A1 _02154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11161__B1 _05223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07904__A1 _02078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11161__C2 _02387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05915__B1 _05767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06183__A3 _00631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10267__A2 _02741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xwrapped_as2650_140 la_data_out[62] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11464__B2 _02028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xwrapped_as2650_151 io_oeb[37] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_182_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_162 la_data_out[53] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XTAP_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10477__I _04376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09409__A1 as2650.stack\[6\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11624_ _03972_ _05663_ _05664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11216__A1 as2650.stack\[10\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06891__A1 _05770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11216__B2 as2650.stack\[9\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11555_ _00773_ _01090_ _04225_ _05601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_129_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08632__A2 _01686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07786__I _02029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06690__I _01132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06643__A1 _00460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10506_ _04583_ _04603_ _04607_ _04618_ _04619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_171_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_144_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11486_ as2650.r123\[3\]\[0\] _05545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_7_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10437_ _02906_ _04549_ _04550_ _04551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_136_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_170_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10368_ _04487_ _04489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_151_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09934__C _03777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_124_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_139_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10299_ _02618_ _02850_ _04434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09506__I net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12038_ _00407_ clknet_leaf_15_wb_clk_i as2650.ins_reg\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_78_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09896__A1 _03774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07026__I _01464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06530_ net5 _00936_ _00974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_111_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07470__B _01902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06865__I _01265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11455__A1 _02089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06461_ _00623_ _00709_ _00903_ _00906_ _00907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_61_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08200_ as2650.stack\[6\]\[11\] _02517_ _02520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_33_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09180_ _03392_ _03400_ _03401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__06882__A1 _01305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06392_ _00476_ _00837_ _00838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_147_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08131_ _02467_ _02468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_147_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09820__A1 _03978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06814__B _01227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06634__A1 _01031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08062_ _02121_ _02415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_88_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07013_ _01308_ _01423_ _01452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_190_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10718__B1 _01828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09584__B1 _03742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06105__I as2650.cycle\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10194__A1 _00778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08964_ as2650.r123_2\[1\]\[7\] _03105_ _03204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08320__I _02627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07915_ _02181_ _02297_ _02269_ _02300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_4719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08895_ _03133_ _03137_ _03139_ _03140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_44_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07846_ _02053_ _02227_ _02246_ _02047_ _00057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_151_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09639__A1 _03797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07777_ _02188_ _02189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_71_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11446__A1 _01889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06775__I _01216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06728_ _05745_ _05782_ _05783_ _05708_ _01171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_140_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09516_ _00648_ _02593_ _03680_ _03681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_71_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11446__B2 as2650.r123\[2\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08311__A1 _02610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__10297__I _03877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09447_ _02534_ _03621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_164_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06659_ _00955_ _01103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08862__A2 _01112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_146_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06873__A1 _01234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09378_ _03568_ _03562_ _03569_ _03570_ _00265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_55_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08329_ _02513_ _02628_ _02633_ _02635_ _00151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_71_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08614__A2 _01501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09811__A1 _00822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06625__A1 _01061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11340_ as2650.stack\[1\]\[7\] _05257_ _05223_ as2650.stack\[3\]\[7\] as2650.stack\[2\]\[7\]
+ _02387_ _05432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_192_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_153_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11271_ as2650.stack\[4\]\[5\] _05210_ _05364_ _05365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_106_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08378__A1 _02663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10222_ _04337_ _04359_ _04371_ _03786_ _00308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_10_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06015__I _00473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10185__A1 _02893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10185__B2 _00507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07050__A1 _01485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10153_ _02586_ _04303_ _04304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_160_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08230__I _02534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10084_ _02212_ _04008_ _04236_ _04237_ _04238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_48_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10488__A2 _04582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08386__B _02671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11437__A1 _01721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11437__B2 as2650.r123\[2\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10986_ _00805_ _05084_ _05085_ _05086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_188_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08853__A2 _00745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06864__A1 _01001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11607_ _05579_ _04444_ _05649_ _05650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_141_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06616__A1 net50 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10412__A2 _03598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_1918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11538_ _05556_ _05578_ _05585_ _04298_ _05586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_116_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06092__A2 _00550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11469_ _00884_ _04349_ _05062_ _05529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_7_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07041__A1 _01432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07465__B _01872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07592__A2 _01104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input9_I io_in[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05961_ _05814_ _05734_ _00420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_24_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09869__A1 _01465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07700_ _05687_ _02121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_78_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10479__A2 _03821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08680_ _02932_ _02952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_38_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_61_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05892_ as2650.r123\[2\]\[6\] as2650.r123_2\[2\]\[6\] _05713_ _05746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_96_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07631_ _01203_ _02042_ _02058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_54_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07562_ _01768_ _01990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_94_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09097__A2 _01648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11745__CLK clknet_4_8_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09301_ _03040_ _03508_ _03510_ _03511_ _00247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06513_ _00956_ _00957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_34_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10100__A1 _03789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07493_ _01920_ _01921_ _01924_ _01925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_62_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_61_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09232_ _03449_ _03450_ _03451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_194_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_146_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06444_ _00822_ _00858_ _00889_ _00890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_181_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10651__A2 _04755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09163_ _03365_ _03367_ _03384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06375_ _00472_ _00819_ _00820_ _00446_ _00821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__11895__CLK clknet_leaf_96_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06607__A1 _01001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08114_ as2650.stack\[0\]\[4\] _02440_ _02455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10403__A2 _03712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09094_ _01546_ _01651_ _03317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_148_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07280__A1 _01605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08045_ _02077_ _02402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_162_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10167__A1 _00891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07032__A1 _01459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09996_ _04150_ _04151_ _04152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_5217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07583__A2 _01080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06386__A3 _00767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08050__I _02256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08947_ _01501_ _03178_ _03188_ _03189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_4505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08878_ _03121_ _03123_ _03124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_56_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07829_ net71 _02235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_3859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07886__A3 _02034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10840_ _02193_ _04914_ _04945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11419__A1 as2650.stack\[9\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10890__A2 _04993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07099__A1 _01393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10771_ _04877_ _04878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_18_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08599__A1 net79 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_193_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_176_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_165_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_165_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11323_ _04409_ _01693_ _00914_ _05415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_154_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_141_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11254_ _05281_ _05348_ _00363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_101_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10158__A1 _00631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09012__A2 _00826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10205_ _00580_ _04347_ _04338_ _04355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__09563__A3 _00816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11185_ _00696_ _05281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_122_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10136_ _04270_ _04103_ _04104_ net92 _01291_ _04288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__06782__B1 _01222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10067_ _04218_ _04220_ _04145_ _04221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__11768__CLK clknet_leaf_92_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08523__A1 as2650.stack\[9\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08523__B2 as2650.stack\[8\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10330__A1 _00737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07877__A3 _02254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_32_wb_clk_i_I clknet_4_7_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06629__B _01072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10881__A2 _04976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07304__I _01739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_189_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10969_ _05055_ _04228_ _02331_ _05070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_56_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06160_ _00586_ _00604_ _00618_ _00619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_156_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_12_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_156_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07262__A1 _01697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06065__A2 _00484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06091_ as2650.cycle\[1\] _00550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_195_1759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09003__A2 _02495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_158_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07014__A1 _01451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09850_ _00698_ _04009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_98_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09554__A3 _03700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10333__C _04458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08762__A1 as2650.stack\[1\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_71_wb_clk_i_I clknet_4_11_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08801_ _03047_ _03041_ _03048_ _03049_ _00209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_140_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09781_ _03888_ _03940_ _03941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06993_ _01432_ _01433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_171_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05944_ _05791_ _05793_ _05798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_6_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08732_ _02692_ _02995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08514__A1 _01733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08663_ _02930_ _01611_ _02931_ _02932_ _02934_ _02935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_26_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05875_ _05724_ _05728_ _05729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_38_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07614_ _02040_ _02042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10872__A2 _04102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08594_ _02866_ _02867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06540__A3 _00983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07545_ _01598_ _01975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08817__A2 _00982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10085__B1 _04238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06828__A1 _00426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07476_ _01888_ _01720_ _01908_ _00025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_22_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10624__A2 _01815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08293__A3 _00495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09215_ _03377_ _03405_ _03430_ _03433_ _03434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_06427_ _00851_ _00872_ _00845_ _00873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_104_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09146_ _03365_ _03367_ _03368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__09778__B1 _03842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06358_ _00805_ _00801_ _00646_ _00806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_120_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08045__I _02077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_194_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09077_ _01626_ _01657_ _03299_ _03300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_139_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06289_ as2650.cycle\[7\] _00691_ _00742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_49_wb_clk_i clknet_4_13_0_wb_clk_i clknet_leaf_49_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_08028_ _02387_ _02388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_155_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11337__B1 _05157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_77_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08753__A1 _02097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_5036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_162_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09979_ _00719_ _04130_ _04134_ _03995_ _03777_ _04135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_39_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output48_I net48 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11941_ _00310_ clknet_leaf_56_wb_clk_i as2650.addr_buff\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_4379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_176_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11872_ _00241_ clknet_leaf_41_wb_clk_i as2650.r123_2\[2\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10823_ _00627_ _05721_ _04929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08808__A2 _03054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_116_wb_clk_i_I clknet_4_2_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06819__A1 _01254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10615__A2 _04722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10754_ _04025_ _03744_ _04862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_125_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09481__A2 _03647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07492__A1 _01784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10685_ _01291_ _04794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_40_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11040__A2 _01111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08992__A1 as2650.stack\[7\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11306_ as2650.stack\[2\]\[6\] _05156_ _05257_ as2650.stack\[1\]\[6\] _05399_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_153_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11237_ as2650.stack\[2\]\[4\] _05296_ _05297_ as2650.stack\[0\]\[4\] _05174_ _05332_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_84_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07547__A2 _01974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08744__A1 as2650.stack\[1\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11168_ _05151_ _05265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_67_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10551__A1 _04590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10119_ _04255_ _04118_ _04120_ _04202_ _04271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_42_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11099_ _02813_ _05190_ _05196_ _05197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_62_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_5581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09514__I _03653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_36_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07180__B1 _01591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_147_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07330_ _01765_ _01766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_16_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10606__A2 _04711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_182_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07261_ _05796_ _01147_ _01698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07483__A1 as2650.stack\[5\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09000_ as2650.stack\[7\]\[4\] _03228_ _03225_ _03235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06212_ _00662_ _00670_ _00671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_121_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_176_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07192_ _01555_ _01557_ _01629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_157_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_1512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06038__A2 _00496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06143_ _00601_ _05702_ _00602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__11031__A2 _00872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_1556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06074_ _00532_ _00533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11933__CLK clknet_leaf_61_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09902_ _00896_ _04043_ _04059_ _04060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_132_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09527__A3 _00581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07538__A2 _01859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09833_ _02612_ _03850_ _03991_ _03992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_141_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09852__C _04010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06210__A2 _00663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09764_ _00704_ _03925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06976_ _01398_ _01416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_27_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08715_ as2650.stack\[15\]\[3\] _02972_ _02983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05927_ _05780_ _05781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__11098__A2 _01204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09695_ _03836_ _03856_ _03857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_26_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05858_ _05711_ _05712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08646_ as2650.stack\[9\]\[7\] _02913_ _02795_ as2650.stack\[8\]\[7\] as2650.stack\[11\]\[7\]
+ _02799_ _02918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XPHY_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07710__A2 _02092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08577_ _02849_ _02850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_145_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_35_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10058__B1 _04211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07879__I _02269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_161_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07528_ as2650.r123\[0\]\[6\] _01958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_167_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09463__A2 _03620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07459_ as2650.stack\[6\]\[11\] _01855_ _01856_ as2650.stack\[4\]\[11\] _01892_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_155_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10470_ _00800_ _04583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09215__A2 _03405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06029__A2 _00448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09129_ _03327_ _03329_ _03351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__11022__A2 _04379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08974__A1 _01686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_155_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10781__A1 _04875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_190_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11022_ _00864_ _04379_ _05121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08726__A1 as2650.stack\[15\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10533__A1 _02057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06201__A2 _00650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08378__C _02671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11924_ _00293_ clknet_leaf_49_wb_clk_i net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10836__A2 _04469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11855_ _00002_ clknet_leaf_47_wb_clk_i as2650.cycle\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_33_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11806__CLK clknet_leaf_134_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07789__I _02200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08394__B _02682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06693__I _01135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10806_ _04875_ _04789_ _04910_ _04911_ _04912_ _00351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_158_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11786_ _00169_ clknet_leaf_85_wb_clk_i as2650.stack\[2\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09454__A2 _02536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06268__A2 _00720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08662__B1 _02933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10737_ _04844_ _04845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11261__A2 _04837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_186_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11104__I _00774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10668_ as2650.stack\[3\]\[4\] _01738_ _01786_ _04778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_12_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11013__A2 _00979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10599_ _03921_ _03920_ _04710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_103_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08965__A1 _05796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07768__A2 _02178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_182_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08717__A1 _02402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08717__B2 _02984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10524__A1 _01845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06728__B1 _05783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08193__A2 _02514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09390__A1 _03542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06830_ _01271_ _01272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__09390__B2 _03580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09244__I _03446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07940__A2 _02297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06761_ _01201_ _01204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_95_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05951__A1 _05760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08500_ _02341_ _02566_ _02772_ _02337_ _02773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_110_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06692_ _01134_ _01135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09480_ _03646_ _02759_ _03647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10827__A2 _04915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08431_ _02710_ _02711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_63_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08362_ _02651_ _02659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_36_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07313_ _01741_ _01729_ _01749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__06259__A2 _00632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08293_ _00735_ _00490_ _00495_ _00501_ _02593_ _02602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
XANTENNA__11252__A2 _05330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_192_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10058__C _04004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_192_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07244_ _01676_ _01680_ _01681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_109_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07175_ _01602_ _01145_ _01606_ _01612_ _01027_ _01613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__11004__A2 _00657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_175_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08956__A1 _02835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06126_ _00544_ _00585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_195_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_156_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_191_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_172_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06057_ _00514_ _00515_ _00516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_47_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05883__S _05736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10515__A1 as2650.stack\[3\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10515__B2 as2650.stack\[2\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09381__A1 _02129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09816_ net35 _03975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_28_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11617__C _00756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07931__A2 _02220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09747_ _03906_ _03907_ _03908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_60_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06959_ _01344_ _01389_ _01398_ _01399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__05942__A1 _05730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11829__CLK clknet_4_7_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10818__A2 _04921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09678_ _03730_ _03791_ _03839_ _03840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_3_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09684__A2 _03845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06498__A2 _00941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08629_ _02823_ _02901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_15_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07695__A1 _01598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11640_ _00023_ clknet_leaf_36_wb_clk_i as2650.r123\[0\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08239__A3 _02547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07447__A1 _01784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11571_ _02956_ _04416_ _05617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11243__A2 _05266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_10_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08942__B _03072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_64_wb_clk_i clknet_4_14_0_wb_clk_i clknet_leaf_64_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__06018__I _05684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10522_ as2650.stack\[13\]\[1\] _01829_ _01826_ as2650.stack\[12\]\[1\] _04635_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_195_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10453_ _00520_ _04566_ _04567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05857__I _05710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06462__B _05677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_170_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08947__A1 _01501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10384_ _04489_ _04500_ _04502_ _00339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_108_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10754__A1 _04025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06422__A2 _00677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11594__I _02956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08389__B _02671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09372__A1 as2650.stack\[3\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11005_ _02607_ _00598_ _05103_ _05104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_42_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07922__A2 _02178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09124__A1 _03305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07686__A1 _02107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11907_ _00276_ clknet_leaf_69_wb_clk_i as2650.ivec\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_146_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_181_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11838_ _00221_ clknet_leaf_105_wb_clk_i as2650.stack\[7\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_76_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_159_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11769_ _00152_ clknet_leaf_92_wb_clk_i as2650.stack\[4\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_159_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06110__A1 _00568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06661__A2 _00835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_155_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_127_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_157_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06949__B1 _01342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10745__A1 _04025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06413__A2 _00844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08980_ _02143_ _02438_ _03218_ _03219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__07982__I _02350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07931_ _02304_ _02220_ _02310_ _02306_ _00078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_68_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10622__B _02907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09363__A1 as2650.stack\[3\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06598__I _01041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07862_ as2650.stack\[12\]\[9\] _02258_ _02259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_84_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11170__A1 as2650.stack\[13\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09601_ _03763_ _01019_ _03740_ _03765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_111_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07913__A2 _02292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11170__B2 as2650.stack\[15\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06813_ _00430_ _05808_ _05792_ _01255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_2
XFILLER_68_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07793_ net87 _02204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09115__A1 _05697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09532_ _05697_ _00840_ _00870_ _02555_ _03696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_83_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06744_ _01176_ _01175_ _01187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__07126__B1 _01563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08469__A3 _00855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06675_ _00429_ _05809_ _01118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_24_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09463_ as2650.stack\[5\]\[6\] _03620_ _03632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08414_ _02675_ _02690_ _02694_ _02698_ _00173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_12_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09394_ _03550_ _03575_ _03581_ _03583_ _00268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_71_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11225__A2 _01445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08345_ _02645_ _02646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_142_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10433__B1 _01744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08276_ _00659_ _01723_ _02550_ _02585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__06101__A1 _00458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10984__A1 _02235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07227_ _01663_ _01664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_180_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11528__A3 _05571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_180_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07158_ _01592_ _01594_ _01595_ _01596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_106_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_145_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10736__A1 _02116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06109_ net7 _00568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_156_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06404__A2 _00849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07601__A1 _02027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07089_ _01506_ _01509_ _01527_ _01528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_160_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11651__CLK clknet_leaf_134_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_4_4_0_wb_clk_i_I clknet_3_2_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_111_wb_clk_i clknet_4_3_0_wb_clk_i clknet_leaf_111_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_82_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11161__A1 as2650.stack\[5\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11161__B2 as2650.stack\[7\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05915__A1 _05766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05915__B2 _05718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output30_I net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12007__CLK clknet_4_2_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09612__I _00632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_130 la_data_out[43] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__11464__A2 _04415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xwrapped_as2650_141 io_oeb[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_128_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_147_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_152 la_data_out[32] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XTAP_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_163 la_data_out[55] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_31_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10672__B1 _01779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06340__A1 _00781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09409__A2 _03577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_145_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11623_ _02616_ _04448_ _04449_ _05661_ _05663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_19_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06891__A2 _00664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11216__A2 _05268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_129_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10424__B1 _02794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11554_ _02756_ _02731_ _05600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_183_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10505_ _04609_ _04582_ _04617_ _04333_ _04618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__10493__I _04374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07840__A1 _02239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11485_ _01772_ _05541_ _05544_ _05540_ _00727_ _00398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_155_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09059__I _01954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10436_ as2650.stack\[13\]\[0\] _01789_ _01793_ as2650.stack\[12\]\[0\] _04550_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__10727__A1 _01844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09593__A1 _02745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10367_ _04481_ _04486_ _04488_ _04405_ _00336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10298_ _01262_ _04432_ _04433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_97_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12037_ _00406_ clknet_leaf_51_wb_clk_i as2650.r123\[3\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11257__C _03813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06159__A1 _00507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07356__B1 _01791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09896__A2 _04053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_187_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11455__A2 _00866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06460_ _00905_ _00906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_178_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06882__A2 _01315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08608__B1 _02876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06391_ _05685_ _00837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07977__I _02345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08130_ _02466_ _02467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_175_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10966__A1 _00444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09820__A2 _01428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08061_ _02412_ _02406_ _02413_ _02414_ _00104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_88_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07012_ _05802_ _01451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_134_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_161_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10718__A1 as2650.stack\[2\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_192_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10718__B2 as2650.stack\[1\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09584__A1 _03740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09584__B2 _03732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06398__A1 _00590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10194__A2 _02008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11391__A1 _02680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08963_ _03191_ _03203_ _00217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_97_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09336__A1 _03044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07914_ as2650.stack\[10\]\[6\] _02293_ _02299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_4709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08894_ _03138_ _03112_ _03087_ _03139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11143__A1 _00775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07347__B1 _01761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09887__A2 _04040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07347__C2 _01782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06121__I _00579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07845_ as2650.stack\[13\]\[12\] _02242_ _02246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07898__A1 _02051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07776_ _02187_ _02188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__05960__I _05752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09432__I _01975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09515_ _00865_ _00787_ _03678_ _03679_ _03680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_37_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06727_ _01169_ _00655_ _01170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11446__A2 _05499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08311__A2 _02614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_1773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09446_ _03614_ _03620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06658_ _01101_ _01102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_1784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08862__A3 _03108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09377_ _03239_ _02653_ _03543_ _03570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06589_ _01027_ _01032_ _01033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_142_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07887__I _02277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08328_ as2650.stack\[4\]\[9\] _02634_ _02635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__11630__C _00712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08614__A3 _01589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08259_ _02567_ _02568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_181_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11202__I _05159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11270_ _05159_ _05364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_180_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10709__A1 _02351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08378__A2 _02667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10221_ _03977_ _04359_ _04370_ _04371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_101_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10185__A2 _04325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11382__A1 _02672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output78_I net78 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10152_ _02549_ _02578_ _03696_ _04303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_133_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10262__B _04301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09327__A1 as2650.stack\[4\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10083_ _00800_ _04237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_134_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09878__A2 _01473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_181_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05870__I _05723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06561__A1 _00722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07063__S _00968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11437__A2 _05499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10985_ _00804_ _05079_ _05085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_16_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08853__A3 _01024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06864__A2 _00966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07797__I _02187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11606_ _05638_ _04443_ _05649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08066__A1 _01770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10948__A1 _04333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11697__CLK clknet_leaf_123_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_195_1908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07813__A1 _02189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11537_ _05579_ _05580_ _05584_ _05585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06616__A2 net78 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11112__I _01914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06206__I _00664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11468_ _02578_ _04353_ _05528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_158_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_193_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09566__A1 _02037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10419_ _04532_ _04533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_174_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11399_ _02003_ _02146_ _02438_ _05475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_135_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_61_wb_clk_i_I clknet_4_14_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07041__A2 _00830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09318__A1 _03020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09318__B2 _03524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05960_ _05752_ _05814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09869__A2 _01457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05891_ _05718_ _05745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_17_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07630_ _02056_ _02057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_53_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07561_ _01988_ _01989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_98_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09300_ as2650.stack\[2\]\[4\] _03504_ _03500_ _03511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_62_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06512_ _00645_ _00558_ _00956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_146_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07492_ _01784_ _01922_ _01923_ _01924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_80_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09231_ _03390_ _03425_ _03450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_107_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06855__A2 _01296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06443_ _00659_ _00861_ _00877_ _00888_ _00889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_179_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_194_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09162_ _03349_ _03366_ _03383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_147_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06374_ _00474_ _00745_ _00820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_9_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08057__A1 _02409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07104__I0 as2650.r123\[0\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07500__I as2650.r123\[0\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_30_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08113_ _02423_ _02454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06607__A2 _01050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09093_ _03314_ _03315_ _03316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_135_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10403__A3 _03705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08044_ _02399_ _02386_ _02400_ _02401_ _00100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_190_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05955__I _05784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10167__A2 _04317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_115_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07032__A2 _01137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09995_ _04137_ _04147_ _04149_ _04151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_88_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_142_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09309__A1 as2650.stack\[2\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07583__A3 _05787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06386__A4 _00831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08946_ _03178_ _03187_ _03188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_88_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11116__A1 _05209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06791__A1 _00423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08877_ _01161_ _03122_ _03123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07828_ _02233_ _02234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__06786__I _01067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11419__A2 _05478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07759_ _02174_ _02156_ _02164_ _02175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_25_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10627__B1 _02795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_183_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_106_wb_clk_i_I clknet_4_3_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10770_ _04875_ _04876_ _04877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_164_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09429_ _03607_ _00279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_55_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06310__A4 _00760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08048__A1 _02402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07410__I _01844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06454__C _05678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09796__A1 _00717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08599__A2 _01671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11322_ _05238_ _01696_ _05414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07271__A2 _01707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06026__I _00484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09765__C _03925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05901__S0 _05705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_180_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09548__A1 _00703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10771__I _04877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11253_ _03279_ _05125_ _05347_ _05348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_122_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05865__I _05718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10704__C _04418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10204_ _03688_ _03714_ _03704_ _04353_ _04354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XANTENNA__08220__A1 _02505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11184_ _03974_ _05280_ _00361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_121_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10135_ _04279_ _04286_ _04287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_121_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06782__A1 as2650.r123\[1\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11107__A1 _02745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06782__B2 _01223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10066_ _00633_ _04219_ _04220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_134_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08397__B _02682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_188_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09720__A1 _03860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08523__A2 _02785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06696__I _01138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10330__A2 _02845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_91_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10618__B1 _01752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10968_ _05061_ _05063_ _05068_ _05069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_62_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09800__I _00688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10094__A1 net41 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11551__B _01038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_147_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10899_ _05001_ _05002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_148_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08039__A1 as2650.stack\[12\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09236__B1 _03454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10167__B _03598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07320__I _01755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_1705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10397__A2 _04511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_145_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06090_ _00548_ _00549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_172_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07262__A2 _00934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_1749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06470__B1 _00915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09539__A1 _00901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10681__I _03661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11346__A1 as2650.stack\[12\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08211__A1 as2650.stack\[6\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_154_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08800_ _02461_ _02475_ _03021_ _03049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_140_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08762__A2 _03004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09780_ _02858_ _01429_ _03939_ _03940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XTAP_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06992_ _05741_ _01432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_136_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08731_ _02415_ _02985_ _02993_ _02994_ _00194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_152_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05943_ _05749_ _05797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_26_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_22_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08662_ _01992_ _01310_ _02933_ _02610_ _02934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_96_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_66_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05874_ _05727_ _05728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06525__A1 _00944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07613_ _02040_ _02041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_93_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08593_ _00880_ _02865_ _02866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_82_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11862__CLK clknet_leaf_27_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07544_ _01964_ _01967_ _01973_ _01883_ _01974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA__08278__A1 _02566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09710__I _03871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10085__A1 _04212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10085__B2 _04161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07475_ _01889_ _01722_ _01853_ _01907_ _01908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_139_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09214_ _03411_ _03408_ _03429_ _03433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_50_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_195_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_194_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06426_ _00871_ _00872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_37_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09778__A1 _02852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09145_ _03349_ _03366_ _03367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_148_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06357_ _00804_ _00805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_108_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09076_ _01628_ _01656_ _03299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_163_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06288_ _00581_ _00740_ _00741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_194_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08027_ _01832_ _02387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11337__A1 as2650.stack\[6\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11337__B2 as2650.stack\[4\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_150_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09950__A1 _04102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08753__A2 _03001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09978_ _04131_ _04133_ _04134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_137_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_18_wb_clk_i clknet_4_5_0_wb_clk_i clknet_leaf_18_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_5059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08929__C _03070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08929_ _03073_ _03170_ _03171_ _03070_ _03172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_4325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07833__C _02201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11940_ _00309_ clknet_leaf_56_wb_clk_i as2650.addr_buff\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11871_ _00240_ clknet_leaf_38_wb_clk_i as2650.r123_2\[2\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_169_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_73_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10822_ _04879_ _04919_ _04924_ _04927_ _04928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_72_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08269__A1 _00734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10076__A1 net87 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06819__A2 _01258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10753_ _00780_ _04859_ _04860_ _04418_ _04861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_129_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10684_ _04792_ _04793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_185_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05893__I3 as2650.r123_2\[0\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11576__A1 _04545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_154_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11305_ as2650.stack\[0\]\[6\] _05297_ _05303_ as2650.stack\[3\]\[6\] _05398_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_181_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11591__A4 _05634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11328__A1 _02592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11735__CLK clknet_leaf_108_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11236_ as2650.stack\[1\]\[4\] _05162_ _05163_ as2650.stack\[3\]\[4\] _05331_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_122_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09941__A1 _04078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08744__A2 _03004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11167_ _00755_ _05264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10551__A2 _04661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10118_ as2650.addr_buff\[4\] _04270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_67_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11098_ _05129_ _01204_ _05195_ _02819_ _05196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_27_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10049_ _04124_ _04126_ _04202_ _04203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_48_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07180__A1 _01565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07180__B2 _01299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_51_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07260_ _00793_ _01697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07483__A2 _01914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_108_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06211_ _00500_ _00669_ _00670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07191_ _01539_ _01560_ _01627_ _01628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__05884__I3 as2650.r123_2\[0\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11567__A1 _01327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06142_ _00480_ _00601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_157_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08432__A1 _02663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10625__B _02907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06073_ _00530_ as2650.cycle\[2\] _00531_ _00532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_160_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11319__A1 _03609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09901_ _04025_ _03872_ _00817_ _04041_ _03925_ _04059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_160_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09832_ _03760_ _03991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09932__A1 _04087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_140_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09705__I _03866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09763_ _02855_ _00683_ _03742_ _03886_ _03924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_86_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06975_ _01086_ _01413_ _01414_ _01088_ _01415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_100_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_4_9_0_wb_clk_i_I clknet_3_4_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12131__I net85 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08714_ _02399_ _02970_ _02981_ _02982_ _00189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_73_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05926_ as2650.r0\[1\] _05780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09694_ _03819_ net93 _03856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09696__B1 _03857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08645_ _02915_ _02916_ _01844_ _02917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_82_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05857_ _05710_ _05711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_55_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08576_ _02848_ _02849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_26_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__12040__CLK clknet_leaf_9_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09440__I _03614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07527_ _01931_ _01910_ _01957_ _00027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_145_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10058__B2 _03995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09999__A1 _03873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11191__B _05192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07474__A2 _01904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07458_ as2650.stack\[7\]\[11\] _01858_ _01859_ as2650.stack\[5\]\[11\] _01891_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_50_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06409_ _05701_ _00767_ _00855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_195_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07389_ _01823_ _01824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_148_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07895__I _02277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09128_ _01644_ _03349_ _03350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_135_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11758__CLK clknet_leaf_80_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08423__A1 as2650.stack\[1\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10535__B _02070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10230__A1 _02806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09059_ _01954_ _03285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_124_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10781__A2 _00628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06304__I _00754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09923__A1 _04078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11021_ _03646_ _04309_ _05119_ _00959_ _05120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08726__A2 _02978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output60_I net60 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10533__A2 _04531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09615__I _00730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_131_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09151__A2 _03372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11923_ _00292_ clknet_4_6_0_wb_clk_i net24 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_45_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11854_ _00001_ clknet_leaf_54_wb_clk_i as2650.cycle\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10049__A1 _04124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10805_ _00711_ _04912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06907__C _01165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10496__I _04608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11246__B1 _05178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11785_ _00168_ clknet_leaf_84_wb_clk_i as2650.stack\[2\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_57_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10736_ _02116_ _04843_ _04844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__06268__A3 _00722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08662__A1 _01992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07465__A2 _01858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08662__B2 _02610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_161_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10667_ as2650.stack\[1\]\[4\] _01814_ _01817_ as2650.stack\[0\]\[4\] as2650.stack\[2\]\[4\]
+ _01875_ _04777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_142_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08414__A1 _02675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09611__B1 _03772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10598_ _04708_ _04709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_154_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10221__A1 _03977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08717__A2 _02970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11219_ _05265_ _05314_ _05315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_190_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06728__A1 _05745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06728__B2 _05708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09390__A2 _03575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11276__B _05369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06760_ _01136_ _01203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_5390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05951__A2 _05727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09142__A2 _03363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06691_ _05781_ _01134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_188_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07153__A1 _01461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08430_ _02709_ _02710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_64_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_145_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11237__B1 _05297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08361_ _02645_ _02658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_75_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07312_ as2650.stack\[7\]\[8\] _01740_ _01747_ as2650.stack\[6\]\[8\] _01748_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_08292_ _00912_ _02595_ _02598_ _02600_ _00753_ _02601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_20_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08653__A1 _02805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11900__CLK clknet_leaf_73_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_1589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07243_ _01576_ _01583_ _00825_ _01679_ _01680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__10460__A1 _03723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08405__A1 _01770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07174_ _01611_ _01147_ _01144_ _01612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_118_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10212__A1 _03647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06125_ _00556_ _00567_ _00572_ _00583_ _00584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_118_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11030__I _05103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06056_ _00454_ _00515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_105_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06431__A3 _00875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09905__A1 _04023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10515__A2 _01835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09815_ _00727_ _03974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09381__A2 _02653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09746_ _02081_ _01310_ _03907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06958_ _01397_ _01398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_100_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10279__A1 _01022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05909_ _05760_ _05734_ _05761_ _05719_ _05762_ _05739_ _05763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XTAP_2005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09677_ _02055_ _01141_ _03839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_2016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06889_ _01267_ _00989_ _01329_ _00654_ _01330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__07144__A1 _01480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08628_ _02882_ _02899_ _02884_ _02900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_2049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08892__A1 _01297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_168_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08559_ _02813_ _02816_ _02817_ _02831_ _02832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XTAP_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_52_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11570_ _05612_ _05613_ _05615_ _00839_ _05616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08644__A1 as2650.stack\[2\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_180_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08942__C _03183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10521_ as2650.stack\[15\]\[1\] _01810_ _01823_ as2650.stack\[14\]\[1\] _04634_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_122_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10452_ _03745_ _04565_ _04566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_109_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06462__C _00749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10203__A1 _00519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10383_ net46 _04494_ _04501_ _04502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_163_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_163_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_33_wb_clk_i clknet_4_7_0_wb_clk_i clknet_leaf_33_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_151_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06422__A3 _00763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_137_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11164__C1 _05223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09345__I _03543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11004_ _03243_ _00657_ _05103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_133_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11906_ _00275_ clknet_leaf_69_wb_clk_i as2650.ivec\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11923__CLK clknet_4_6_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10690__A1 _04397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11837_ _00220_ clknet_leaf_104_wb_clk_i as2650.stack\[7\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_61_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11768_ _00151_ clknet_leaf_92_wb_clk_i as2650.stack\[4\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_92_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10442__A1 _04076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10719_ _04540_ _04826_ _04827_ _04828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__10954__I net69 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11699_ _00082_ clknet_leaf_123_wb_clk_i as2650.stack\[10\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06110__A2 as2650.last_intr vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10993__A2 _05090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06661__A3 _01104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09060__A1 _03285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10745__A2 _04009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06949__B2 _01333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_170_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07930_ as2650.stack\[11\]\[11\] _02307_ _02310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_114_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07861_ _02250_ _02258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__05909__C1 _05762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09600_ _03740_ _03763_ _01018_ _03764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_116_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11170__A2 _05266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06812_ _01252_ _01123_ _01253_ _01254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_110_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07792_ _02189_ _02197_ _02201_ _02203_ _00046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_37_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09531_ _00832_ _02567_ _02738_ _03694_ _00778_ _03695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XANTENNA__11458__B1 _05513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06743_ _01185_ _01068_ _01070_ _01186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_42_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07126__A1 as2650.r123\[1\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07931__C _02306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08469__A4 _02741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09462_ _03565_ _03627_ _03630_ _03631_ _00288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06674_ _00999_ _01099_ _01113_ _01117_ _00014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__08874__A1 _01139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_51_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07503__I _01824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08413_ as2650.stack\[1\]\[10\] _02697_ _02698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_51_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09393_ _02364_ _03579_ _03582_ _03583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_36_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08344_ _02644_ _02645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_178_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10433__A1 as2650.stack\[11\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10433__B2 as2650.stack\[10\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08275_ _00860_ _02583_ _02584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_149_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06101__A2 _00557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_177_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10984__A2 _00808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07226_ _05724_ _01663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_138_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09426__I0 as2650.ivec\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_193_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_175_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_4_1_0_wb_clk_i clknet_3_0_0_wb_clk_i clknet_4_1_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_49_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07157_ _01565_ _01017_ _01595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09874__B _04031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_156_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_118_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06108_ _00560_ _00566_ _00567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_195_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07088_ _01520_ _01526_ _01527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__07601__A2 _02028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06039_ _00497_ _00498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_121_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07365__A1 _01105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11161__A2 _05257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11946__CLK clknet_leaf_54_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09729_ _03842_ _03843_ _03889_ _03890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_47_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xwrapped_as2650_120 io_out[33] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06325__C1 _00690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xwrapped_as2650_131 la_data_out[45] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_70_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output23_I net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_142 io_oeb[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_167_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xwrapped_as2650_153 la_data_out[34] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XANTENNA__10672__A1 as2650.stack\[15\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_164 la_data_out[57] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XANTENNA__10672__B2 as2650.stack\[14\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06340__A2 _00789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11622_ net85 _05661_ _05662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_42_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10424__A1 as2650.stack\[5\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11553_ _05108_ _05598_ _05599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_11_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10424__B2 as2650.stack\[4\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09290__A1 _02368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_195_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10504_ _04610_ _04615_ _04616_ _04617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_109_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07840__A2 _02207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11484_ _02028_ _05543_ _05544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_137_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10435_ as2650.stack\[15\]\[0\] _04536_ _04542_ as2650.stack\[14\]\[0\] _04549_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_183_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09593__A2 _00748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10366_ net43 _04487_ _04488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_154_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_51_wb_clk_i_I clknet_4_13_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06699__I _01141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10297_ _03877_ _04432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_97_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09075__I _03297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12036_ _00405_ clknet_leaf_57_wb_clk_i as2650.r123\[3\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_120_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07356__A1 as2650.stack\[14\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07356__B2 as2650.stack\[13\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11455__A3 _00657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_181_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06390_ _00511_ _00835_ _00836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_21_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08608__B2 _02879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_193_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06619__B1 _05778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10415__A1 _04305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_187_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10684__I _04792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08084__A2 _02427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11720__D _00103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_90_wb_clk_i_I clknet_4_8_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_147_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08060_ _02181_ _02258_ _02385_ _02414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_179_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07011_ _01388_ _01450_ _00018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_146_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09033__A1 _01847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10718__A2 _04542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09584__A2 _00683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06398__A2 _05702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10194__A3 _04343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11391__A2 _05467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08962_ _01563_ _03177_ _03202_ _03099_ _03203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_142_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08103__B _02446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07913_ _02102_ _02292_ _02296_ _02298_ _00072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__09336__A2 _03533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08893_ _01034_ _03138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_111_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11143__A2 _01249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07347__B2 as2650.stack\[8\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07942__B _02316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07844_ _02239_ _02220_ _02245_ _02241_ _00056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_84_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07775_ _02186_ _02031_ _02034_ _02187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_56_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09514_ _03653_ _03679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_25_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06726_ as2650.holding_reg\[1\] _01169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__08847__A1 _03092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09445_ _02284_ _02541_ _03619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06657_ _01100_ _01101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_129_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_185_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09376_ as2650.stack\[3\]\[6\] _03552_ _03569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06588_ _01028_ _01029_ _01031_ _01032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_127_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08327_ _02626_ _02634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09272__A1 _01975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08075__A2 _02425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06086__A1 _00543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08258_ _00557_ _02004_ _02567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06625__A3 _01068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07209_ as2650.r0\[1\] _01542_ _01646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_10_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09024__A1 _03098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08189_ _02511_ _02512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_152_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10709__A2 _04792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10220_ _00707_ _00736_ _04360_ _04369_ _04370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_3_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07586__A1 _01080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11382__A2 _05457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10151_ _03721_ _04300_ _04302_ _00306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_79_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_192_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_160_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09327__A2 _03521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10082_ _04235_ _04236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_82_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_135_wb_clk_i_I clknet_4_1_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10342__B1 _04458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06010__A1 _00467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10893__A1 _03662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10893__B2 _04996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06561__A2 _01004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10984_ _02235_ _00808_ _05084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_28_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10645__A1 _03958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_31_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06982__I _01421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06864__A3 _01128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09498__C _00697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11605_ _00824_ _02903_ _02860_ _05647_ _05648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_30_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09263__A1 _02345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08066__A2 _02249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11536_ _04626_ _05565_ _05583_ _02621_ _05566_ _05584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__07813__A2 _02220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10009__I _02893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09015__A1 _00848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11467_ _00702_ _05526_ _02581_ _05527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_87_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09566__A2 _01041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10418_ _04469_ _03757_ _04532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_136_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11549__B _04501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11398_ _02151_ _05467_ _05474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07577__A1 _00554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10349_ _00670_ _03673_ _02741_ _04472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_124_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10581__B1 _02913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06222__I _00679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_140_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12019_ _00388_ clknet_leaf_105_wb_clk_i as2650.stack\[9\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_39_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05890_ _05743_ _05727_ _05744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_39_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_54_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06552__A2 _00987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07560_ _01987_ _01988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_94_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08829__A1 _00744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06511_ _05714_ _00955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10636__A1 net58 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07491_ as2650.stack\[15\]\[12\] _01874_ _01900_ as2650.stack\[13\]\[12\] _01923_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_94_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07988__I _02199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09230_ _03414_ _03448_ _03449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_146_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06442_ _00882_ _00883_ _00660_ _00887_ _00888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_167_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09161_ _03352_ _03370_ _03381_ _03382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_166_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11641__CLK clknet_leaf_36_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06373_ _00512_ _00816_ _00818_ _00819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__08057__A2 _02406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07104__I1 as2650.r123_2\[0\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08112_ _02402_ _02436_ _02451_ _02453_ _00116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__07002__B _01013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07265__B1 _01699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09092_ _03312_ _03313_ _03315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_120_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08043_ _02167_ _02392_ _02397_ _02401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_174_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_147_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09708__I _00638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07568__A1 _01985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09994_ _04147_ _04149_ _04137_ _04150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_103_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09309__A2 _03504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08945_ _03186_ _01458_ _03125_ _03187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_135_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08517__B1 _01751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08876_ _03062_ _03122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_111_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07827_ _01543_ _02233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06543__A2 _00554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07740__A1 _01984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07758_ _02096_ _02174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_53_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06709_ _01139_ _01140_ _01149_ _01151_ _00943_ _01152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__10627__A1 as2650.stack\[13\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10627__B2 as2650.stack\[12\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07689_ _02102_ _02092_ _02103_ _02111_ _00035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_38_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09428_ as2650.ivec\[4\] _03279_ _03604_ _03607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_158_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09359_ as2650.stack\[3\]\[2\] _03546_ _03556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06059__A1 _00513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06307__I _00685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11321_ _00756_ _05413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_177_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_107_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05901__S1 _05753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09618__I _03781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09548__A2 _01712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08522__I _02794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11252_ _00757_ _05330_ _05337_ _05346_ _05278_ _05347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_153_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07559__A1 _00605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10203_ _00519_ _03713_ _02759_ _04349_ _04353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_155_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11183_ _03267_ _05125_ _05279_ _05280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_161_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10134_ _04004_ _04285_ _03781_ _04286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_7_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_5731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11107__A2 _04651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06782__A2 _01116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10065_ _04217_ _04214_ _04215_ _04219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10618__A1 as2650.stack\[7\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10618__B2 as2650.stack\[5\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09484__A1 _02732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08287__A2 _00481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10967_ _04802_ _05056_ _05065_ _05067_ _02350_ _05068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__11664__CLK clknet_leaf_121_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06298__A1 _00747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10898_ _02217_ _05000_ _05001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_31_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09236__B2 _03107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11123__I _00823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09787__A2 _03946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07798__A1 as2650.stack\[14\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_1717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11519_ _02777_ _05560_ _05567_ _05568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_144_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09528__I _02017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06470__A1 _00508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09539__A2 _02004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06470__B2 _00891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11346__A2 _02271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06991_ _01297_ _01431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07970__A1 _02332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08730_ as2650.stack\[15\]\[7\] _02978_ _02969_ _02994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__06887__I _05766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05942_ _05730_ _05795_ _05796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_132_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08661_ net1 _02933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__10857__A1 _04157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05873_ _05726_ _05727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_82_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07612_ _02021_ _02040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_93_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08592_ _02722_ _02865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_35_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07543_ _01968_ _01969_ _01972_ _01973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_41_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08278__A2 _02569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06836__B _00944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11282__A1 _05298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07474_ _01890_ _01904_ _01906_ _01849_ _01907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_22_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07511__I _01791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09213_ _03162_ _03298_ _03432_ _00238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06425_ _00666_ _00871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_167_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09144_ _05742_ _01360_ _03366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11034__A1 _02028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_194_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09778__A2 _01302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06127__I _00585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06356_ _00601_ _00804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_147_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11585__A2 _05625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09075_ _03297_ _03298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06287_ _00518_ _00681_ _00740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_30_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_190_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09438__I _03612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06461__A1 _00623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08026_ _02385_ _02386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_146_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11337__A2 _05212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10545__B1 _04653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_89_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09950__A2 _04089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09977_ _04132_ _04088_ _04133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_104_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07961__A1 _02329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08928_ _01445_ _03074_ _03171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_4315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10848__A1 _04175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08859_ as2650.r123_2\[1\]\[0\] _03105_ _03106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_185_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11870_ _00239_ clknet_leaf_38_wb_clk_i as2650.r123_2\[2\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10821_ _04725_ _04925_ _04926_ _04927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_72_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_183_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09466__A1 _02184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08269__A2 _01037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10752_ _04811_ _04844_ _04860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11273__A1 as2650.stack\[2\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06819__A3 _01260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08674__C1 _01460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07421__I _01746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10683_ _04007_ _04791_ _04792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_71_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06037__I _00495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11576__A2 _04552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06452__A1 _00589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11304_ _05209_ _05395_ _05396_ _05397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_4_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11235_ _05813_ _05282_ _05321_ _05329_ _05330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_101_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09941__A2 _04097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11166_ _05259_ _05262_ _05222_ _05263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_136_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07952__A1 _02323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10117_ _03721_ _04268_ _04269_ _00305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_95_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_4_14_0_wb_clk_i clknet_3_7_0_wb_clk_i clknet_4_14_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_5550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11097_ _05129_ _05194_ _05195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10839__A1 _04913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10048_ as2650.addr_buff\[0\] _04173_ as2650.addr_buff\[2\] _04202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__06500__I _00943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11118__I _05215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08901__B1 _03130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07180__A2 _01011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11562__B _02752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09457__A1 _03509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10957__I _05057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11999_ _00368_ clknet_4_15_0_wb_clk_i as2650.r123_2\[3\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_90_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07468__B1 _01879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10178__B _04328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06210_ _05704_ _00663_ _05694_ _00668_ _00669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XANTENNA__11016__A1 _00880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07190_ _01540_ _01559_ _01627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_121_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09686__C _00533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06141_ _00508_ _00599_ _00600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_117_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07487__B _01846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08432__A2 _02707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_172_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06072_ net6 _00531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_195_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11319__A2 _05189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09900_ _00810_ _04056_ _04057_ _03917_ _04058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_144_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09831_ _03987_ _03988_ _03989_ _03990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_119_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06974_ _01392_ _01412_ _01414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09762_ _03734_ _03920_ _03922_ _03923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_58_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08111__B _02446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07506__I _01827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05925_ _05776_ _05725_ _05777_ _05717_ _05778_ _05706_ _05779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
X_08713_ _02449_ _02974_ _02979_ _02982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09693_ _03848_ _03854_ _03855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09696__A1 _03793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08644_ as2650.stack\[2\]\[7\] _02909_ _01733_ _02916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_2209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05856_ _05709_ _05710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_55_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09721__I _03718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08575_ _01271_ _02848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10867__I _04469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09448__A1 as2650.stack\[5\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_81_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07526_ _01932_ _01911_ _01853_ _01956_ _01957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__11255__A1 _04129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10058__A2 _04208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07459__B1 _01856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09999__A2 _04134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08120__A1 _02409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07457_ _01726_ _01890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06408_ _00848_ _00850_ _00853_ _00854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__11007__A1 _02568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07388_ _01822_ _01823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_195_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11558__A2 _05603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09127_ _05731_ _01510_ _03349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06339_ _00451_ _00789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_178_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09620__A1 _03723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08423__A2 _02689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_105_wb_clk_i clknet_4_3_0_wb_clk_i clknet_leaf_105_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_157_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_194_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09058_ _03271_ _03284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10230__A2 _02747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08072__I _02423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08009_ _02200_ _02373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_191_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10518__B1 _01826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08187__A1 _02198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11020_ _03646_ _00904_ _02349_ _05119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_89_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09923__A2 _03850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07934__A1 as2650.stack\[11\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output53_I net94 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11922_ _00291_ clknet_leaf_49_wb_clk_i net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_4189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10777__I _04877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11382__B _05461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11853_ _00013_ clknet_4_12_0_wb_clk_i as2650.cycle\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09439__A1 _02003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10049__A2 _04126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11246__A1 as2650.stack\[10\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10804_ as2650.ivec\[2\] _04470_ _04841_ _04878_ _04873_ _04911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_11784_ _00167_ clknet_leaf_85_wb_clk_i as2650.stack\[2\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11246__B2 as2650.stack\[9\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08111__A1 _02452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10735_ _04007_ _04791_ _04843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_158_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08662__A2 _01310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_185_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06673__A1 as2650.r123\[1\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06990__I _01393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10666_ _01764_ _04774_ _04775_ _04776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__11702__CLK clknet_leaf_116_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09611__A1 _03759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10597_ _03750_ _04708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08414__A2 _02690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10221__A2 _04359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_181_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11218_ _05309_ _05313_ _05314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_9_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11182__B1 _05263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06728__A2 _05782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10524__A3 _04636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_1_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11149_ _02135_ _05245_ _05135_ _05246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_95_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07326__I _01752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06230__I _00687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11485__A1 _01772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06690_ _01132_ _01133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_97_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08360_ _02519_ _02646_ _02652_ _02657_ _00160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__11237__A1 as2650.stack\[2\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11237__B2 as2650.stack\[0\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07311_ _01746_ _01747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_3_wb_clk_i clknet_4_1_0_wb_clk_i clknet_leaf_3_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_60_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08291_ _00506_ _02599_ _02597_ _02600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_32_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08653__A2 _02924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07242_ _01572_ _01678_ _01679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_137_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10460__A2 _04570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07929__C _02306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07173_ _01610_ _01611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_88_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08405__A2 _02138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06124_ _00573_ _00582_ _00583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10212__A2 _00700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06967__A2 _01236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_172_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06055_ _05720_ _00514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_132_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08620__I _00677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11173__B1 _05269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06719__A2 _01161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07916__A1 _02113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09814_ _03971_ _03973_ _00298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_86_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09118__B1 _03340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09745_ _02080_ net11 _03906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06957_ _01392_ _01396_ _01397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_112_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05908_ as2650.r123\[1\]\[4\] as2650.r123\[0\]\[4\] as2650.r123_2\[1\]\[4\] as2650.r123_2\[0\]\[4\]
+ _05683_ _05736_ _05762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XANTENNA__10279__A2 _03877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11476__A1 _00729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06888_ _05727_ _00988_ _01328_ _01329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09676_ net89 net10 _03838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_95_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_54_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08341__A1 as2650.stack\[4\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08627_ _01182_ _01407_ _02876_ _02898_ _02899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_05839_ _05692_ _05693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10597__I _03750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08892__A2 _03113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11228__A1 _00955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08067__I _02418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08558_ _02819_ _02825_ _02830_ _02831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_74_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11725__CLK clknet_leaf_86_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07509_ _01739_ _01940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_51_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08489_ _00754_ _02761_ _02762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_167_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07447__A3 _01880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08644__A2 _02909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10520_ _04626_ _04631_ _04632_ _04633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_161_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10451__A2 _00687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_167_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10451_ _03739_ _00687_ _04565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_10_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10382_ _00678_ _04501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_184_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_41_wb_clk_i_I clknet_4_6_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07080__A1 _01020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09626__I _00552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07907__A1 as2650.stack\[10\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11164__B1 _02271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11003_ _00864_ _03648_ _03686_ _05101_ _05102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_46_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11808__D _00191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11164__C2 as2650.stack\[3\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_73_wb_clk_i clknet_4_10_0_wb_clk_i clknet_leaf_73_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_120_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08686__B _02351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11467__A1 _00702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07590__B _02017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08332__A1 _02516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11905_ _00274_ clknet_leaf_72_wb_clk_i as2650.stack\[6\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_185_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11219__A1 _05265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10690__A2 _00895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11836_ _00219_ clknet_leaf_104_wb_clk_i as2650.stack\[7\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11767_ _00150_ clknet_leaf_92_wb_clk_i as2650.stack\[4\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_80_wb_clk_i_I clknet_4_10_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10442__A2 _03731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10718_ as2650.stack\[2\]\[5\] _04542_ _01828_ as2650.stack\[1\]\[5\] _04827_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_11698_ _00081_ clknet_leaf_123_wb_clk_i as2650.stack\[11\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06110__A3 net75 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10649_ _04394_ _00896_ _04725_ _04758_ _04759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_155_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08399__A1 as2650.stack\[2\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06225__I _00682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06949__A2 _01239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_100_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10903__C _04419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09899__A1 _04041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11155__B1 _05248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07860_ _02197_ _02252_ _02253_ _02257_ _00060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__05909__B1 _05761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05909__C2 _05739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06811_ _01015_ _00432_ _01227_ _01253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_56_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07791_ as2650.stack\[14\]\[8\] _02202_ _02203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_68_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11458__A1 _01707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06742_ _01072_ _01185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09530_ _00878_ _00490_ _00669_ _02550_ _03694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_37_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07126__A2 _01116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08323__A1 _02138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_188_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09461_ _02110_ _02536_ _03612_ _03631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06673_ as2650.r123\[1\]\[0\] _01116_ _01117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_97_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06885__A1 _00437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08412_ _02688_ _02697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_145_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09392_ _02511_ _03582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_24_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08343_ _02249_ _02630_ _02644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09823__A1 _01466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11898__CLK clknet_leaf_72_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06637__A1 _01080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08274_ _00863_ _02582_ _02583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10433__A2 _04536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07225_ _01660_ _01661_ _01662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_140_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09426__I1 _03273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_192_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07156_ _01319_ _01593_ _01594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_161_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10197__A1 _00548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06107_ _00563_ _00565_ _00566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07062__A1 _01096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07087_ _01523_ _01524_ _01525_ _01526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__07675__B _02063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_160_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10813__C _04651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09446__I _03614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06038_ _05676_ _00496_ _00497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_105_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08350__I _02650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_125_wb_clk_i_I clknet_4_0_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07989_ _02356_ _02357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09728_ _01273_ _01254_ _01258_ _01260_ _03889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_41_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08314__A1 _02606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xwrapped_as2650_110 io_oeb[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_09659_ _00629_ _03821_ _03822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xwrapped_as2650_121 io_out[34] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__06325__C2 _00775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_132 la_data_out[47] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_82_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xwrapped_as2650_143 io_oeb[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_128_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06876__A1 _01316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_154 la_data_out[36] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_82_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05923__I0 as2650.r123\[2\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xwrapped_as2650_165 la_data_out[59] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_42_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output16_I net16 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11621_ _02340_ _05660_ _05661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_168_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xclkbuf_leaf_120_wb_clk_i clknet_4_2_0_wb_clk_i clknet_leaf_120_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_30_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06628__A1 _01015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11621__A1 _02340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10424__A2 _02784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11552_ _03657_ _01498_ _02748_ _05598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_36_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10276__B _04412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09290__A2 _03502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_184_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10503_ _02846_ _04586_ _04616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11483_ _05264_ _05542_ _03780_ _05543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_155_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10434_ _04540_ _04546_ _04547_ _04548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_137_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10188__A1 _00563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07053__A1 _00500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10727__A3 _04835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10365_ _04480_ _04487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_163_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06800__A1 _01180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08260__I _02568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10296_ _04426_ _04430_ _04431_ _00322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_156_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_191_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12035_ _00404_ clknet_leaf_53_wb_clk_i as2650.r123\[3\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_2_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07356__A2 _01746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10360__A1 _00881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_150_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10112__A1 _04109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11455__A4 _03100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10663__A2 _04760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05914__I0 as2650.r123\[1\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_178_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11819_ _00202_ clknet_leaf_107_wb_clk_i as2650.stack\[1\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09805__A1 _00629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06619__A1 _05720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_186_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06619__B2 _05708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11612__A1 _02805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10186__B _04336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06095__A2 as2650.cycle\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07010_ _01225_ _01449_ _01450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_174_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_162_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10179__A1 net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10914__B _04570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07044__A1 _05740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08792__A1 as2650.stack\[8\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08961_ _01589_ _03178_ _03201_ _03202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_69_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07912_ _02177_ _02297_ _02269_ _02298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08892_ _01297_ _03113_ _03135_ _03136_ _03137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_96_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08544__A1 _01462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07347__A2 _01762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07843_ as2650.stack\[13\]\[11\] _02242_ _02245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_112_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10351__A1 _00697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07774_ _02132_ _02186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_42_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09513_ _02823_ _02568_ _03678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_25_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06725_ _00434_ _01167_ _01168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_37_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11036__I _00847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10654__A2 _05761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09444_ _03542_ _03613_ _03616_ _03618_ _00283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06656_ _01022_ _01100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_168_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06587_ net50 _01030_ _01031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_52_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09375_ _02112_ _03568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_178_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_181_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08326_ _02505_ _02628_ _02629_ _02633_ _00150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__08345__I _02645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11603__A1 _02737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_166_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09272__A2 _02234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_177_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06086__A2 _00544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08257_ _00506_ _02566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_53_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07208_ _01635_ _01643_ _01644_ _01645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_153_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08188_ _02510_ _02511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10824__B _00698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_180_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07139_ _01413_ _01400_ _01497_ _01489_ _01577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_106_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08783__A1 as2650.stack\[8\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10150_ net92 _04067_ _04301_ _04302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_106_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11119__B1 _05154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10081_ _03737_ _04227_ _04234_ _03818_ _04235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_173_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09904__I _02745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07338__A2 _01773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10342__A1 _04399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10342__B2 _00827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06010__A2 _00468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10893__A2 _04975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_16_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10983_ _00622_ _00699_ _05083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_186_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10645__A2 _02955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05879__I _05732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06864__A4 _01304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11604_ _05599_ _05605_ _05644_ _05646_ _05647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_168_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09263__A2 _03465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07274__A1 _01290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11535_ _04462_ _02770_ _05582_ _05583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_128_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09015__A2 _03101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11466_ _00450_ _02768_ _02754_ _02740_ _05526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_183_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_clkbuf_3_3_0_wb_clk_i_I clknet_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10417_ _04530_ _04531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_87_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11397_ _05472_ _05473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_180_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07577__A2 _00904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_152_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10348_ _04406_ _04471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_139_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10581__A1 as2650.stack\[15\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10581__B2 as2650.stack\[13\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10279_ _01022_ _03877_ _04416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12018_ _00387_ clknet_leaf_101_wb_clk_i as2650.stack\[9\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_79_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11565__B _05610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10333__A1 _00737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06552__A3 _00995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08829__A2 _00937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06510_ _00947_ _00953_ _00954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_146_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_146_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07490_ as2650.stack\[14\]\[12\] _01877_ _01879_ as2650.stack\[12\]\[12\] _01922_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__10636__A2 net57 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06441_ _00886_ _00516_ _00887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_94_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_179_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09160_ _03355_ _03369_ _03381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_148_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06372_ _00817_ _00818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_187_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_163_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_148_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08111_ _02452_ _02425_ _02446_ _02453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_159_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06068__A2 _00499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09091_ _03312_ _03313_ _03314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__07265__A1 _01462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08042_ as2650.stack\[12\]\[2\] _02390_ _02400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11936__CLK clknet_leaf_61_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07937__C _02158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07017__A1 _01454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_176_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07509__I _01739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07568__A2 _01989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09993_ _03932_ _03963_ _04148_ _04149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__10572__A1 _01787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_192_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08944_ _03184_ _03185_ _03186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_48_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08517__A1 as2650.stack\[3\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08517__B2 as2650.stack\[1\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_4519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08875_ _01136_ _03111_ _03072_ _03120_ _03121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_111_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07826_ _02222_ _02231_ _02232_ _02201_ _00051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_84_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11194__C _05241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06543__A3 _00986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07757_ as2650.stack\[11\]\[4\] _02149_ _02173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_44_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06708_ _01150_ _01046_ _01040_ _01151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__10627__A2 _01751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07688_ _02104_ _02110_ _01997_ _02111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_52_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09493__A2 _03643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08296__A3 _02604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09427_ _03606_ _00278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06639_ _01061_ _01062_ _01068_ _01083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_25_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09358_ _02066_ _03555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_166_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06059__A2 _00517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08309_ _02331_ _02618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_138_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_176_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09289_ _02665_ _03502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_142_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11320_ _05281_ _05412_ _00365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_10_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_165_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10554__B _04374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11251_ _05264_ _05345_ _05346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09548__A3 _02580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08756__A1 as2650.stack\[1\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07559__A2 _00974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10202_ _03710_ _03697_ _04346_ _04351_ _04352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_136_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06323__I _00773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11182_ _00757_ _05255_ _05263_ _05277_ _05278_ _05279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_192_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_106_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10133_ _04283_ _04284_ _04285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_66_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07863__B _02257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09634__I _03796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_125_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10064_ _04214_ _04215_ _04217_ _04218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11385__B _05461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05990__A1 _00448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10866__A2 _04947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11809__CLK clknet_leaf_5_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08694__B _02965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06993__I _01432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10618__A2 _01839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10966_ _00444_ _05066_ _05067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09484__A2 _03650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06298__A2 _05678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11291__A2 _01589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10897_ _04222_ _04974_ _05000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_182_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11959__CLK clknet_4_5_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09236__A2 _03340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07247__A1 _01059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07247__B2 _01092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_156_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07798__A2 _02208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11518_ _02571_ _05564_ _05565_ _02780_ _05566_ _05567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_89_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06470__A2 _00599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11449_ _05503_ _05513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08747__A1 _02449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07329__I _01764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10554__A1 _04432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_193_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06990_ _01393_ _01430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input7_I io_in[35] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07970__A2 _00853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05941_ _05741_ _05749_ _05786_ _05794_ _05795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_113_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05981__A1 _05813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10306__A1 _01905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05872_ _05725_ _05726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__10857__A2 _04930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08660_ _00792_ _02932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_66_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06525__A3 _00968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07611_ _02038_ _02039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_26_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08591_ _02809_ _02840_ _02843_ _02863_ _02864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_81_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06930__B1 _01370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07999__I _02200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07542_ _01766_ _01970_ _01971_ _01972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_34_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07473_ _01905_ _01803_ _01906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_179_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_161_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09212_ as2650.r123_2\[2\]\[3\] _03342_ _03431_ _03107_ _03432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__10358__C _04479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_182_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06424_ _00505_ _00834_ _00870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_56_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_194_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09143_ as2650.r0\[7\] _01218_ _03365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06355_ _00671_ _00802_ _00770_ _00803_ _00007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_33_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08986__A1 as2650.stack\[7\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09074_ _00514_ _03067_ _03297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_175_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06286_ _00711_ _00739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10374__B _04301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08025_ _02255_ _02385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_162_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06461__A2 _00709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11189__C _03859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10545__A1 _00446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_143_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_5006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09976_ net37 _04132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_130_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07961__A2 _02279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08927_ _01430_ _03111_ _03169_ _03170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_131_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11636__D _00019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05972__A1 _05771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09163__A1 _03365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08858_ _03104_ _03105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08910__A1 _03149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07809_ _02217_ _02218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_29_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08789_ _02090_ _03040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_2925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10820_ _04157_ _04102_ _04926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_96_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09466__A2 _03617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08674__B1 _01138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10751_ _04023_ _03733_ _04858_ _04859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11273__A2 _05225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_98_wb_clk_i clknet_4_9_0_wb_clk_i clknet_leaf_98_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__08674__C2 _01435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10320__I1 as2650.holding_reg\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_27_wb_clk_i clknet_4_7_0_wb_clk_i clknet_leaf_27_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__06318__I _00768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10682_ net60 _04746_ _04791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__07229__A1 _01029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_142_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08533__I _00878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06988__B1 _01425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10284__B _00765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_154_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11303_ as2650.stack\[5\]\[6\] _05302_ _05303_ as2650.stack\[7\]\[6\] _05396_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_154_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08729__A1 _02381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11234_ _03815_ _05327_ _05328_ _05329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06053__I _00511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10536__A1 _04646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11165_ _05216_ _05260_ _05261_ _05262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_68_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10731__C _00732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10116_ _04256_ _04067_ _04165_ _04269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_49_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11096_ _01725_ _04638_ _05193_ _05194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_5540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09154__A1 _03129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11631__CLK clknet_leaf_37_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10047_ _04175_ _04176_ _04201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__10303__I _02855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10839__A2 _04531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08901__A1 _01222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08901__B2 as2650.r123_2\[1\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08708__I _02971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11998_ _00367_ clknet_leaf_52_wb_clk_i as2650.r123_2\[3\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11781__CLK clknet_leaf_85_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09457__A2 _03617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10949_ _05035_ _05050_ _04948_ _05051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_127_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09209__A2 _03428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06140__A1 _00496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_176_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07768__B _02140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06140_ _00496_ _00598_ _00599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_8_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_157_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10775__A1 _02125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06071_ as2650.cycle\[10\] _00530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06443__A2 _00861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07059__I _01088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09393__A1 _02364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09830_ _03987_ _03988_ _03849_ _03989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_28_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_150_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09761_ _03886_ _03921_ _03922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06973_ _01392_ _01412_ _01413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_132_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08712_ as2650.stack\[15\]\[2\] _02972_ _02981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05924_ as2650.r123\[1\]\[0\] as2650.r123\[0\]\[0\] as2650.r123_2\[1\]\[0\] as2650.r123_2\[0\]\[0\]
+ as2650.ins_reg\[0\] _05711_ _05778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XANTENNA__10213__I _00702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09692_ _03850_ _03852_ _03853_ _03854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09696__A2 _03855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08643_ as2650.stack\[1\]\[7\] _02913_ _02914_ as2650.stack\[0\]\[7\] as2650.stack\[3\]\[7\]
+ _02799_ _02915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_05855_ net51 _05709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_167_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_184_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08574_ _02846_ _02847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_82_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09448__A2 _03620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_35_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07525_ _01890_ _01953_ _01955_ _01802_ _01956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__07459__A1 as2650.stack\[6\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11255__A2 _01474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08656__B1 _01436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08120__A2 _02454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07456_ _01351_ _01889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_126_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06407_ _00852_ _00853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_22_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11007__A2 _02731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07387_ _01779_ _01822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08959__A1 _01596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09126_ _03316_ _03332_ _03347_ _03348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06338_ _00781_ _00783_ _00787_ _00788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_104_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08353__I _02644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_175_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09620__A2 _03725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10766__A1 as2650.ivec\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10766__B2 _04845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_31_wb_clk_i_I clknet_4_7_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09057_ _03283_ _00231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06269_ _00711_ _00719_ _00723_ _00724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_108_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07631__A1 _01203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08008_ _02078_ _02357_ _02371_ _02372_ _00093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_117_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10518__A1 as2650.stack\[9\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_191_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10518__B2 as2650.stack\[8\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11654__CLK clknet_leaf_3_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08187__A2 _02491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06198__A1 _05680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11191__A1 _02000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10551__C _02334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07934__A2 _02160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09959_ _04068_ _04114_ _04115_ _00301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__05945__A1 _05735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_8_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10123__I _03991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output46_I net46 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09912__I _03724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07698__A1 _02104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11921_ _00290_ clknet_leaf_97_wb_clk_i as2650.stack\[5\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_185_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07860__C _02257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_174_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11852_ _00012_ clknet_leaf_67_wb_clk_i as2650.cycle\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_61_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07432__I _01734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10803_ _04790_ _04878_ _04909_ _00732_ _04910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__11246__A2 _05225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11783_ _00166_ clknet_leaf_85_wb_clk_i as2650.stack\[2\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_186_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08111__A2 _02425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_70_wb_clk_i_I clknet_4_11_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10734_ _02107_ _04789_ _04840_ _04842_ _00739_ _00349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__06122__A1 _00540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06673__A2 _01116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10665_ as2650.stack\[7\]\[4\] _01809_ _01756_ as2650.stack\[4\]\[4\] _04775_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_90_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09611__A2 _03770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10757__A1 _00521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10596_ _00446_ _04703_ _04706_ _04604_ _04707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_166_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08178__A2 _02497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_194_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11217_ _05160_ _05311_ _05312_ _05313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_29_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput70 net70 la_data_out[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__10461__C _04363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11182__A1 _00757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06511__I _05714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11148_ _05130_ _05245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_96_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09127__A1 _05731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11079_ _01877_ _05178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_5381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07689__A1 _02102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07689__B2 _02111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11237__A2 _05296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08638__B1 _02909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_4_13_0_wb_clk_i_I clknet_3_6_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07310_ _01745_ _01746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_36_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08290_ _02547_ _02599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06113__A1 _00485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10996__A1 _04532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10996__B2 _03757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07241_ _01461_ _00764_ _01677_ _01678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_108_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07172_ _01609_ _01610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_157_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10748__A1 _04802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_191_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06123_ _00577_ _00580_ _00581_ _00582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_118_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_172_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06054_ _00492_ _00513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_191_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_173_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_28_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_160_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_115_wb_clk_i_I clknet_4_2_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11173__A1 as2650.stack\[14\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11173__B2 as2650.stack\[12\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09813_ _03951_ _03837_ _03972_ _03973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_99_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07916__A2 _02292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10920__A1 _03662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09118__A1 _03108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11039__I _00613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10920__B2 _05022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09744_ _00633_ _03901_ _03904_ _03905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_86_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06956_ as2650.holding_reg\[4\] _00655_ _01395_ _01396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_74_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_189_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05907_ as2650.r123\[2\]\[4\] as2650.r123_2\[2\]\[4\] _05736_ _05761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11483__B _03780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09675_ _03719_ _03837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06887_ _05766_ _01328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_27_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08341__A2 _02627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08626_ _01484_ _01489_ _01074_ _01416_ _02898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_15_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05838_ as2650.alu_op\[1\] _05692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_27_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08557_ _02807_ _01498_ _02829_ _02830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__11228__A2 _05131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10287__I0 _04417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07508_ _01854_ _01935_ _01938_ _01939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__10436__B1 _01793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06104__A1 _00525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08488_ _02758_ _02760_ _02761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_93_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10987__A1 _04400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10987__B2 _00586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06655__A2 _01057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07439_ as2650.stack\[11\]\[10\] _01858_ _01872_ _01873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__07852__A1 _01985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_168_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11502__I _05681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10450_ _04561_ _04562_ _04563_ _04564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08083__I _02423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10739__A1 _04229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09109_ _03319_ _03331_ _03332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__07604__A1 _05675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10381_ _03273_ _04490_ _04499_ _04500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10203__A3 _02759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07080__A2 _01518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09357__A1 _03550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11164__B2 as2650.stack\[0\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11002_ _00725_ _00866_ _03766_ _05101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_105_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07907__A2 _02293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06331__I _00780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10506__A4 _04618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06591__A1 _00609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11393__B _05468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11467__A2 _05526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11904_ _00273_ clknet_leaf_72_wb_clk_i as2650.stack\[6\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07540__B1 _01761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11835_ _00218_ clknet_leaf_32_wb_clk_i as2650.r123_2\[1\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11219__A2 _05314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10427__B1 _01793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08096__A1 as2650.stack\[0\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11766_ _00149_ clknet_leaf_68_wb_clk_i net75 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_158_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_158_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10717_ as2650.stack\[3\]\[5\] _04822_ _01825_ as2650.stack\[0\]\[5\] _04826_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_174_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11697_ _00080_ clknet_leaf_123_wb_clk_i as2650.stack\[11\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_9_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10648_ _04395_ _04587_ _04758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_139_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10579_ _04626_ _04689_ _04690_ _04691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_170_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09817__I _03719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09348__A1 as2650.stack\[3\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11155__A1 _01269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09899__A2 _03820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06241__I _00576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05909__A1 _05760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10902__A1 _04454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06810_ _00430_ _05808_ _05792_ _01252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
X_07790_ _02187_ _02202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06582__A1 _00930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06741_ _01069_ _01073_ _01031_ _01184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_110_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11458__A2 _05502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_168_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09520__A1 _00442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08323__A2 _02630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09460_ as2650.stack\[5\]\[5\] _03615_ _03630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_77_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06672_ _01115_ _01116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_1924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_184_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08411_ _02672_ _02690_ _02694_ _02696_ _00172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_52_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06885__A2 _00656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09391_ as2650.stack\[6\]\[1\] _03577_ _03581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_91_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_181_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08087__A1 _02327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08342_ _02527_ _02639_ _02640_ _02643_ _00156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_127_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_51_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09823__A2 _01458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06637__A2 _00766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08273_ _00992_ _02582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07224_ as2650.holding_reg\[7\] _01486_ _01661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_146_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09587__A1 _03750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07155_ _05797_ _01454_ _01593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_118_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09727__I _03887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_195_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06106_ _00536_ _00564_ _00565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07086_ _05732_ _01109_ _01525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07062__A2 _01480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08631__I _02902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09339__A1 _03047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06037_ _00495_ _00496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08011__A1 _02174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06573__A1 _01016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07988_ _02199_ _02356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_25_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09727_ _03887_ _03888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06939_ _01378_ _01379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_186_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_170_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09511__A1 _00496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08314__A2 _02622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xwrapped_as2650_100 io_oeb[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_09658_ _03729_ _03791_ _03821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
Xwrapped_as2650_111 io_oeb[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__06325__A1 _00623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xwrapped_as2650_122 io_out[35] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__10121__A2 _04124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06325__B2 _00771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08609_ _02872_ _02881_ _02882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xwrapped_as2650_133 la_data_out[48] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xwrapped_as2650_144 io_oeb[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XANTENNA__06876__A2 _01298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09589_ _03749_ _03752_ _03723_ _03753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xwrapped_as2650_155 la_data_out[38] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_128_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_166 la_data_out[61] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XANTENNA__11842__CLK clknet_leaf_102_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06340__A4 _00787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11620_ _04652_ _04399_ _05660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11082__B1 _01962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11551_ _03657_ _05140_ _02768_ _01038_ _05597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__07825__A1 as2650.stack\[14\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_156_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10502_ _00689_ _04613_ _04614_ _04615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_17_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11992__CLK clknet_4_5_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11482_ _04652_ _05522_ _03666_ _05524_ _05542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_155_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10433_ as2650.stack\[11\]\[0\] _04536_ _01744_ as2650.stack\[10\]\[0\] _04547_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_152_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07866__B _02257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10188__A2 _02547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11385__A1 _02675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08541__I _01037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10364_ _01101_ _04483_ _04485_ _04486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08250__A1 _02551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06800__A2 _01188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10295_ as2650.holding_reg\[1\] _04426_ _04431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_78_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11137__A1 _05220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12034_ _00403_ clknet_leaf_57_wb_clk_i as2650.r123\[3\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06061__I _00519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06996__I _01435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10360__A2 _00979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09502__A1 _00825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06316__A1 _05704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05914__I1 as2650.r123\[0\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08069__A1 as2650.stack\[0\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11818_ _00201_ clknet_4_3_0_wb_clk_i as2650.stack\[1\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_72_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06619__A2 _05777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11749_ _00132_ clknet_leaf_88_wb_clk_i as2650.stack\[7\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11612__A2 _04741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10179__A2 _00611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09547__I _03710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07044__A2 _00991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08241__A1 _00992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_192_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08960_ _01619_ _03071_ _03200_ _03127_ _03201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_83_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07911_ _02277_ _02297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_151_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08891_ _02849_ _03059_ _03113_ _03136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_97_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09741__A1 net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08544__A2 _02815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07842_ _02239_ _02214_ _02244_ _02241_ _00055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_151_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08400__B _02682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10351__A2 _04470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07773_ _02122_ _02172_ _02183_ _02185_ _00045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_56_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09512_ _03674_ _03676_ _03677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_37_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06724_ _00664_ _01167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_1710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11300__A1 _02837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07504__B1 _01934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09443_ _02045_ _03617_ _02542_ _03618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06655_ _01000_ _01057_ _01098_ _01099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_164_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_1787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09374_ _03565_ _03562_ _03566_ _03567_ _00264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_52_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06586_ net78 _01030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_33_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08325_ _02632_ _02633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_138_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11603__A2 _02569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__11052__I _05150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06146__I _00459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08256_ _02560_ _02564_ _02565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08480__A1 _00831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_140_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_192_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07207_ as2650.r0\[4\] _01358_ _01644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_137_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10891__I _04622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08187_ _02198_ _02491_ _02471_ _02510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_101_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05985__I _00443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07138_ _01575_ _01576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08361__I _02645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08232__A1 _02521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_161_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_175_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07069_ _01265_ _01200_ _01361_ _01508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_160_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06794__A1 _01234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11119__A1 as2650.stack\[1\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11119__B2 as2650.stack\[3\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10080_ _04209_ _02955_ _04233_ _04234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_47_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09732__A1 _02856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10342__A2 _04463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07705__I _02125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10982_ _02235_ _05081_ _05082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_56_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09920__I _04076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_188_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08536__I _02808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07440__I _01810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11603_ _02737_ _02569_ _05600_ _05645_ _05646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_15_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06056__I _00454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11534_ _05561_ _05578_ _05581_ _05582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_184_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07274__A2 _00848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08471__A1 _02737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09795__C _03789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11465_ _04620_ _05524_ _05221_ _05525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_125_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10734__C _00739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11738__CLK clknet_leaf_114_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08223__A1 _02513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10416_ _04529_ _04530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_178_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11396_ _05459_ _05472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_87_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10030__A1 _03789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09971__A1 _04124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10347_ _04469_ _04470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_139_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10581__A2 _02908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10278_ _02865_ _02844_ _04415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_39_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11888__CLK clknet_leaf_102_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09723__A1 _03836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12017_ _00386_ clknet_leaf_101_wb_clk_i as2650.stack\[9\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_78_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06537__A1 _00973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10333__A2 _04460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10636__A3 net56 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06440_ _00885_ _00886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_62_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_107_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06371_ as2650.addr_buff\[7\] _00575_ _00817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_21_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11597__A1 _05221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08110_ _02086_ _02452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09090_ _05723_ _01212_ _03313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_147_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08462__A1 _00773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06068__A3 _00509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08041_ _02066_ _02399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_147_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10021__A1 _04156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09992_ _03999_ _04138_ _04148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08943_ _01474_ _03063_ _03185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10660__B _04769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08517__A2 _02782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08874_ _01139_ _03112_ _03118_ _03119_ _03120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_130_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06528__A1 _00694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11521__A1 _02618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07825_ as2650.stack\[14\]\[13\] _02188_ _02232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_56_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07756_ _02157_ _02172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_56_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12043__CLK clknet_4_4_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06707_ _00423_ _01150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_44_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07687_ _02109_ _02110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_168_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11922__D _00291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_183_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09426_ as2650.ivec\[3\] _03273_ _03604_ _03606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06638_ _01081_ _01082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_13_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08356__I _02644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06700__A1 _00930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09357_ _03550_ _03544_ _03551_ _03554_ _00260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_55_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_178_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06569_ _01001_ _00981_ _00983_ _01013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__09896__B _03813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11588__A1 _03642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08308_ _02614_ _02616_ _02617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_165_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09288_ _03028_ _03494_ _03499_ _03501_ _00244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_138_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10260__A1 _00639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_193_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08239_ _00524_ _00758_ _02547_ _02548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_140_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07008__A2 _01429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08205__A1 as2650.stack\[6\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08091__I _02435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11250_ _05170_ _05344_ _05345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_120_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_179_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10201_ _04347_ _00740_ _04348_ _04350_ _04351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__06216__B1 _00646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08756__A2 _02998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07559__A3 _01986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09953__B2 _04109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11181_ _05124_ _05278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_133_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10132_ net68 _02940_ _04284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_106_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_5711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_134_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10063_ _04216_ _04217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06519__A1 _00872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07435__I _01791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11512__A1 _00826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05990__A2 _05700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07192__A1 _01555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09650__I _02889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10079__A1 _04228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10965_ _02229_ _05064_ _05066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_44_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_189_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10729__C _04062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06298__A3 _00749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08692__A1 _00865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10896_ _02217_ _04999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_141_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11579__A1 _04652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08444__A1 _02680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10251__A1 _04395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11517_ _02746_ _05566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10237__S _04385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11448_ _01223_ _03454_ _05512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_125_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10003__A1 _03917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08747__A2 _03001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11379_ _02663_ _05457_ _05458_ _05461_ _00375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_158_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10554__A2 _04661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11576__B _05579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05940_ _05741_ _05791_ _05793_ _05749_ _05794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_136_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_117_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11503__A1 _02860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10306__A2 _04439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05981__A2 _00426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07345__I _01780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05871_ _05688_ _05683_ _05725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_15_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07183__A1 _01055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07610_ _02037_ _02038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_66_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08590_ _02842_ _02857_ _02862_ _02863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_38_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06930__A1 as2650.r123\[1\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07541_ as2650.stack\[14\]\[14\] _01782_ _01762_ as2650.stack\[13\]\[14\] _01971_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_81_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_50_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07472_ _01306_ _01905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07486__A2 _01865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11282__A3 _05375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11903__CLK clknet_leaf_72_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09211_ _03410_ _03430_ _03431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__10490__A1 _04584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06423_ _00765_ _00671_ _00768_ _00868_ _00869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_22_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_195_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09142_ _03359_ _03363_ _03364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_148_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08904__I _01234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06354_ _00713_ _00691_ _00803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08435__A1 _02672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10242__A1 _03797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09073_ _03284_ _03295_ _03296_ _00234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_148_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06285_ _00728_ _00738_ _00012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_163_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06997__A1 _01436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08024_ _01983_ _02384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09935__A1 net63 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10545__A2 _04649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09975_ net38 _04131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_103_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_77_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08926_ _01431_ _03133_ _03168_ _03119_ _03169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_4306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05972__A2 _05773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08857_ _00695_ _03099_ _03103_ _03104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XTAP_4339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07174__A1 _01611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07808_ _02216_ _02217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08788_ _03037_ _03022_ _03038_ _03039_ _00206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_57_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07739_ _02151_ _02156_ _02158_ _02159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_44_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08269__A4 _02577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10750_ _01697_ _04056_ _04858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08674__A1 _00626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08674__B2 _01042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10481__A1 _04590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09409_ as2650.stack\[6\]\[6\] _03577_ _03594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_158_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10681_ _03661_ _04790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_90_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07229__A2 _00991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10233__A1 _03655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_67_wb_clk_i clknet_4_12_0_wb_clk_i clknet_leaf_67_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_138_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06988__A1 _01299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10284__C _03749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11302_ as2650.stack\[6\]\[6\] _05156_ _05157_ as2650.stack\[4\]\[6\] _05395_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_142_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11233_ _03149_ _02867_ _03679_ _02860_ _05328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_106_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08729__A2 _02974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07874__B _02264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11164_ as2650.stack\[1\]\[2\] _05257_ _02271_ as2650.stack\[0\]\[2\] _05223_ as2650.stack\[3\]\[2\]
+ _05261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_136_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10115_ _02218_ _03788_ _04267_ _04163_ _04268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_67_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11095_ _02027_ _00874_ _05191_ _05192_ _05193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_5541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05963__A2 _00421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09154__A2 _03298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10046_ _04199_ _04200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_29_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07165__A1 _00928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08901__A2 _03108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11926__CLK clknet_leaf_62_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11997_ _00366_ clknet_leaf_7_wb_clk_i as2650.r0\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_95_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11415__I _05460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10459__C _04225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10948_ _04333_ _05044_ _05049_ _00673_ _05050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__08665__A1 _02342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07468__A2 _01900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10472__A1 _04186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10879_ _04806_ _04982_ _04983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06140__A2 _00598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_118_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10224__A1 _03686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09090__A1 _05723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06979__A1 as2650.holding_reg\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_1516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06070_ _00528_ _00529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09917__A1 _04071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_105_wb_clk_i_I clknet_4_3_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09555__I _03718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10922__C _04912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_193_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09393__A2 _03579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09760_ _01697_ _03921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06972_ _01396_ _01412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08711_ _02394_ _02970_ _02977_ _02980_ _00188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05923_ as2650.r123\[2\]\[0\] as2650.r123_2\[2\]\[0\] _05711_ _05777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09145__A2 _03366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09691_ _01274_ _03849_ _03760_ _03853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__07156__A1 _01319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08642_ _02794_ _02914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05854_ _05707_ _05708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_132_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09504__B _02894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06903__A1 _01342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08573_ _01142_ _02846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_82_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_58_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07524_ _01954_ _01727_ _01955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_63_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06419__I _00864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08656__A1 _02135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07459__A2 _01855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08656__B2 _02927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10463__A1 _04554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07455_ as2650.r123\[0\]\[3\] _01888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_34_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06406_ _00851_ _00657_ _00852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_195_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08408__A1 _02663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07386_ _01766_ _01813_ _01820_ _01821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_124_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09125_ _03319_ _03331_ _03347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05890__A1 _05743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10215__A1 net91 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_194_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08959__A2 _03122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06337_ _00786_ _00787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_175_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09081__A1 _01569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11060__I _05158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10766__A2 _04470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07092__B1 _01530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09056_ _03282_ as2650.r123_2\[0\]\[4\] _03271_ _03283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_136_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_159_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06268_ _00549_ _00720_ _00722_ _00723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_30_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09908__A1 _04041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08007_ _02170_ _02202_ _02366_ _02372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_89_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06199_ _00651_ _00657_ _00658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05993__I _00451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10518__A2 _01829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11176__C1 as2650.stack\[10\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08187__A3 _02471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11191__A2 _00874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09958_ _04087_ _03976_ _02894_ _04115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_103_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05945__A2 _05740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11949__CLK clknet_4_6_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08909_ _03150_ _03151_ _03079_ _03152_ _03153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_135_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09889_ _04046_ _04047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_3402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_114_wb_clk_i clknet_4_2_0_wb_clk_i clknet_leaf_114_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_44_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11920_ _00289_ clknet_leaf_97_wb_clk_i as2650.stack\[5\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_131_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07698__A2 _02119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07713__I _02132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output39_I net39 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11851_ _00011_ clknet_leaf_66_wb_clk_i as2650.cycle\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10802_ _02809_ _04906_ _04908_ _04909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_54_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06329__I _00778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11782_ _00165_ clknet_leaf_88_wb_clk_i as2650.stack\[2\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08647__A1 as2650.stack\[10\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10454__A1 _04156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10733_ as2650.ivec\[0\] _04470_ _04841_ _04793_ _04530_ _04842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_183_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10664_ as2650.stack\[6\]\[4\] _01780_ _01751_ as2650.stack\[5\]\[4\] _04774_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_186_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10206__A1 _03692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05881__A1 _05733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09072__A1 as2650.r123_2\[0\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10595_ _04596_ _04704_ _04705_ _04706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_177_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07083__B1 _01380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_182_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09375__I _02112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11216_ as2650.stack\[10\]\[3\] _05268_ _05178_ as2650.stack\[9\]\[3\] _05312_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_68_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput60 net60 la_data_out[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__07386__A1 _01766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput71 net71 la_data_out[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__11182__A2 _05255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_190_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11147_ _05243_ _04696_ _05244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_172_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_110_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11078_ _05165_ _05177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_5371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_5393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10029_ _03759_ _04180_ _04183_ _03811_ _00552_ _04184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_37_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08886__A1 _03110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11573__C _05140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07689__A2 _02092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07623__I _02049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06239__I _00695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08638__A1 as2650.stack\[7\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08638__B2 as2650.stack\[6\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10445__A1 _04418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_189_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06113__A2 _00571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10996__A2 _05080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07240_ _01568_ _00764_ _01677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08454__I _00602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_192_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07171_ _01608_ _01609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09063__A1 as2650.r123_2\[0\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10748__A2 _04855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06122_ _00540_ as2650.cycle\[12\] _00581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_118_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_195_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06053_ _00511_ _00512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_145_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10652__C _04606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06702__I _01144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11173__A2 _05268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09812_ _02893_ _03972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_154_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09118__A2 _03337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10920__A2 _05002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06955_ _05806_ _00990_ _01394_ _00828_ _01395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_09743_ _03811_ _03903_ _03904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07129__A1 _01565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07961__C _02281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05906_ _05759_ _05760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_100_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09674_ net32 _03836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08877__A1 _01161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06886_ _01077_ _01327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08629__I _02823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08625_ _02896_ _02897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05837_ as2650.alu_op\[2\] _05691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_55_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11055__I _01937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08556_ _02342_ _02826_ _02827_ _02828_ _02829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07507_ as2650.stack\[5\]\[13\] _01936_ _01937_ as2650.stack\[4\]\[13\] _01938_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__10436__A1 as2650.stack\[13\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10287__I1 _01061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10436__B2 as2650.stack\[12\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08487_ _02759_ _01711_ _02760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__11930__D _00299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06104__A2 _00562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10987__A2 _05083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07438_ _01734_ _01872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_10_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05863__A1 as2650.ins_reg\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_195_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07369_ _01728_ _01800_ _01802_ _01804_ _01805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__09054__A1 _03279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10739__A2 _05746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09108_ _03326_ _03330_ _03331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_108_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10380_ _01431_ _04491_ _04499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08801__A1 _03047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07604__A2 _02018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10203__A4 _04349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09039_ _01884_ _03250_ _03268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_124_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08313__B _02621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07708__I _02128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12050_ _00419_ clknet_leaf_18_wb_clk_i net74 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_116_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07368__A1 _01100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11164__A2 _05257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11001_ _00451_ _05098_ _05099_ _00866_ _00754_ _05100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_104_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_191_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06040__A1 _00490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06591__A2 _00947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08539__I _02592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07443__I _01876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11903_ _00272_ clknet_leaf_72_wb_clk_i as2650.stack\[6\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07540__B2 as2650.stack\[12\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11834_ _00217_ clknet_leaf_32_wb_clk_i as2650.r123_2\[1\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_27_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10427__A1 as2650.stack\[1\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10427__B2 as2650.stack\[0\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11765_ _00148_ clknet_leaf_80_wb_clk_i as2650.stack\[5\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_82_wb_clk_i clknet_4_8_0_wb_clk_i clknet_leaf_82_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_18_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08096__A2 _02440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09293__A1 _03033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10978__A2 _05031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10716_ _02906_ _04823_ _04824_ _04825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_92_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11696_ _00079_ clknet_leaf_119_wb_clk_i as2650.stack\[11\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07843__A2 _02242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10647_ _04709_ _04755_ _04756_ _04419_ _04757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_31_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10578_ as2650.stack\[11\]\[2\] _02908_ _04681_ as2650.stack\[10\]\[2\] _04690_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_127_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07618__I _01996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11155__A2 _05241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05909__A2 _05734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10902__A2 _05002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06740_ _00592_ _01175_ _01177_ _01182_ _01082_ _01183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_97_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08449__I _05670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09520__A2 _00782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10666__A1 _01764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06671_ _00695_ _01106_ _01114_ _01115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_36_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08410_ as2650.stack\[1\]\[9\] _02695_ _02696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_58_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09390_ _03542_ _03575_ _03578_ _03580_ _00267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_55_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08341_ as2650.stack\[4\]\[14\] _02627_ _02643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__10418__A1 _04469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_181_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_177_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11644__CLK clknet_leaf_36_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08087__A2 _02430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09284__A1 _03020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10969__A2 _04228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10647__C _04419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08184__I _02506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08272_ _02580_ _02581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_138_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07223_ _01029_ _00871_ _01660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_164_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07154_ _01316_ _01591_ _01592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_121_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09587__A2 _02747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11794__CLK clknet_leaf_86_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07598__A1 as2650.stack\[13\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06105_ as2650.cycle\[4\] _00564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_118_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07085_ _05759_ _01199_ _01524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_195_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07528__I as2650.r123\[0\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06432__I _05704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06036_ _00491_ _00494_ _00495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_47_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09339__A2 _03533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08011__A2 _02202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06022__A1 _00480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07987_ _00728_ _02355_ _00089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__11925__D _00294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06573__A2 _00977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06588__B _01031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07770__A1 as2650.stack\[11\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06938_ as2650.r123\[0\]\[4\] as2650.r123_2\[0\]\[4\] net51 _01378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_09726_ _01002_ _03887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09511__A2 _02548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06869_ net11 _01310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_09657_ _02952_ _03820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_27_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xwrapped_as2650_101 io_oeb[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__06325__A2 _00499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xwrapped_as2650_112 io_oeb[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__10121__A3 _04126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xwrapped_as2650_123 io_out[36] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08608_ _02873_ _02875_ _02876_ _02879_ _02880_ _02881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XTAP_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xwrapped_as2650_134 la_data_out[50] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xwrapped_as2650_145 io_oeb[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_167_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09588_ _03751_ _03752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xwrapped_as2650_156 la_data_out[40] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_187_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10409__A1 _02732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_167 la_data_out[63] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_42_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08539_ _02592_ _02812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08078__A2 _02427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_184_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11082__A1 as2650.stack\[14\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11550_ _02027_ _05588_ _05596_ _00411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_195_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11082__B2 as2650.stack\[15\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_168_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10501_ _04611_ _04612_ _04614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_155_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09027__A1 _05677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11481_ _03977_ _05525_ _05540_ _05541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_183_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09918__I _00626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10432_ as2650.stack\[9\]\[0\] _02784_ _02794_ as2650.stack\[8\]\[0\] _04546_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08822__I _03065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07589__A1 _00470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11385__A2 _05457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10363_ _01139_ _04484_ _04485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_164_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07438__I _01734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06261__A1 _00712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06342__I net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10294_ _04427_ _04429_ _04430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_152_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12033_ _00402_ clknet_leaf_53_wb_clk_i as2650.r123\[3\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_105_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_26_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09653__I _02608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06013__A1 _00459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07761__A1 as2650.stack\[11\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07173__I _01610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10648__A1 _04395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09502__A2 _02352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06316__A2 _00590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_181_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10663__A4 _04772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05914__I2 as2650.r123_2\[1\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08069__A2 _02419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11817_ _00200_ clknet_leaf_107_wb_clk_i as2650.stack\[1\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_57_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_144_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10467__C _04506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11748_ _00131_ clknet_leaf_83_wb_clk_i as2650.stack\[7\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_144_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09018__A1 _01725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10820__A1 _04157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11679_ _00062_ clknet_leaf_131_wb_clk_i as2650.stack\[12\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_179_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11579__B _05610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11376__A2 _02138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08241__A2 _00747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07348__I _01765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_143_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06252__I as2650.cycle\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_142_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07792__B _02201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07910_ as2650.stack\[10\]\[5\] _02293_ _02296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08890_ _00426_ _03134_ _03135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_97_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10887__A1 _03816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07841_ as2650.stack\[13\]\[10\] _02242_ _02244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09741__A2 net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07752__A1 as2650.stack\[11\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07772_ _02184_ _02178_ _02140_ _02185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_22_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06723_ _01165_ _01166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_09511_ _00496_ _02548_ _03675_ _03676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_37_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11300__A2 _05205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07504__B2 as2650.stack\[6\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09442_ _02529_ _03617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_64_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06654_ _01000_ _01097_ _01098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_92_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08907__I _03058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07811__I _02219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09373_ _02110_ _02653_ _03543_ _03567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06585_ _05730_ _01029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_33_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08324_ _02631_ _02632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_142_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_193_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09009__A1 as2650.stack\[7\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08255_ _02561_ _02563_ _02564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_165_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08480__A2 _00768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06871__B _01144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07206_ as2650.r0\[5\] _01216_ _01643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_101_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08186_ as2650.stack\[6\]\[8\] _02507_ _02509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08642__I _02794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07137_ _01573_ _01574_ _01575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_165_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06243__A1 _00520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07068_ _01328_ _01200_ _01361_ _01507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__11001__C _00754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11119__A2 _05153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06794__A2 _00829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06019_ _00476_ _00477_ _00478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_153_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07743__A1 _02060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09709_ _03870_ _03743_ _03871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10981_ _04595_ _05078_ _05067_ _05081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09496__A1 _02809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_output21_I net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07721__I _02140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09248__A1 _01597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11602_ _02764_ _02740_ _03638_ _05633_ _05645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_93_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06337__I _00786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10802__A1 _02809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11533_ _01262_ _05522_ _05192_ _02350_ _05581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__07274__A3 _01104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08471__A2 _02569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06482__A1 _00529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11464_ _05520_ _04415_ _05521_ _02028_ _05523_ _05524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_109_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10415_ _04305_ _04519_ _04528_ _04529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_87_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11395_ _02686_ _05467_ _05468_ _05471_ _00381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_152_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10566__B1 _04675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06072__I net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10346_ _03692_ _04469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_151_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09971__A2 _04126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_171_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10277_ _01008_ _04412_ _04414_ _04405_ _00320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_97_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09383__I _02510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12016_ _00385_ clknet_leaf_101_wb_clk_i as2650.stack\[9\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09723__A2 _03837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10869__A1 _04167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06537__A2 _00975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_4_0_0_wb_clk_i clknet_3_0_0_wb_clk_i clknet_4_0_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_53_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10097__A2 _04229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10636__A4 net55 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11153__I _01219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11046__A1 _00760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06370_ _00815_ _00816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_148_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_175_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11597__A2 _04696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_147_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08462__A2 _00964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06068__A4 _00526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09558__I _02037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08040_ _02394_ _02386_ _02395_ _02398_ _00099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_163_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09411__A1 _03568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_192_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10021__A2 _04124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09991_ _04046_ _04139_ _04147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_157_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11832__CLK clknet_leaf_27_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08942_ _01954_ _03111_ _03072_ _03183_ _03184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_142_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout88_I net64 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08411__B _02694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10660__C _04588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08873_ _03057_ _03119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_97_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06528__A2 _00971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07725__A1 _01991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07824_ _02230_ _02231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_84_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09478__A1 _00564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07755_ _02078_ _02141_ _02169_ _02171_ _00041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_37_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06706_ _01142_ _00934_ _01145_ _01148_ _01149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_53_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11285__A1 _05152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08637__I _01822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07686_ _02107_ _02083_ _02108_ _02109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_129_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08150__A1 _02325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_50_wb_clk_i_I clknet_4_13_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06637_ _01080_ _00766_ _01081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_25_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09425_ _03605_ _00277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_164_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11063__I _01870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06157__I _00615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06568_ _00427_ _01011_ _01012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09356_ as2650.stack\[3\]\[1\] _03552_ _03553_ _03554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_21_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11588__A2 _04462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08307_ _02615_ _02616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09287_ as2650.stack\[2\]\[1\] _03496_ _03500_ _03501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06499_ _00935_ _00939_ _00942_ _00943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_20_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05996__I _00447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08238_ _00992_ _00734_ _02547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_20_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10260__A2 _04392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08372__I _02665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_153_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08169_ _02487_ _02497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_146_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10200_ _00548_ as2650.cycle\[7\] _00525_ _04349_ _04350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__06216__A1 _00462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11180_ _05264_ _05276_ _05277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_190_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10131_ _04215_ _04280_ _04282_ _04283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_106_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output69_I net69 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06620__I _00988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10062_ net66 _01608_ _04216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_88_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_102_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07716__A1 _02135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10079__A2 _04232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10964_ _02229_ _05064_ _05065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_28_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08141__A1 _02318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_182_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_188_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08692__A2 _02807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10895_ _04223_ _04700_ _04997_ _04998_ _04912_ _00354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_31_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11028__A1 _04409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11705__CLK clknet_leaf_114_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05900__S _05753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11579__A2 _02614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_145_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09641__A1 _01041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08444__A2 _02717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_184_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06455__A1 _00862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10251__A2 _04392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_106_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11516_ _03641_ _05243_ _02570_ _05565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_195_1709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11447_ _05510_ _05511_ _00393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_109_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11378_ _05460_ _05461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_125_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07955__A1 _02325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10329_ _04456_ _04458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07707__A1 _01980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11503__A2 _00751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05870_ _05723_ _05724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11267__A1 _02613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07540_ as2650.stack\[15\]\[14\] _01832_ _01761_ as2650.stack\[12\]\[14\] _01970_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08457__I _00948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08132__A1 as2650.stack\[8\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07471_ _01893_ _01896_ _01903_ _01883_ _01904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_165_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_195_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09210_ _03411_ _03429_ _03430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_06422_ _00865_ _00677_ _00763_ _00867_ _00868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_22_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09141_ _03361_ _03362_ _03363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_37_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_134_wb_clk_i_I clknet_4_1_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06353_ _00781_ _00801_ _00802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08435__A2 _02707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06446__A1 _00891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09072_ as2650.r123_2\[0\]\[7\] _03259_ _03296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10242__A2 _04387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08192__I _02506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06284_ _00468_ _00570_ _00733_ _00737_ _00738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_135_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08023_ _02122_ _02373_ _02382_ _02383_ _00097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_190_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_163_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10227__I _03750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06461__A4 _00906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09935__A2 net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10671__B _01786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07946__A1 _02318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09974_ _04024_ _04122_ _04128_ _04129_ _04130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08141__B _02474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10950__B1 _05033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12010__CLK clknet_leaf_117_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06440__I _00885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08925_ _01599_ _03113_ _03167_ _03078_ _03168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_170_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09699__A1 _02070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11058__I _01942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05972__A3 _00430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08856_ _03102_ _03103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_111_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08371__A1 _02186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07807_ net67 _02216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_85_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05999_ _00457_ _00458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08787_ _02452_ _02475_ _03031_ _03039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_2905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11258__A1 net52 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07738_ _02157_ _02158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11728__CLK clknet_leaf_115_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08123__A1 _02461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08674__A2 _01601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07669_ net60 _02093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_53_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06685__A1 _00637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09408_ _03565_ _03589_ _03592_ _03593_ _00272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_80_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10481__A2 _04592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10680_ _04530_ _04789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_129_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11878__CLK clknet_leaf_99_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09339_ _03047_ _03533_ _03538_ _03539_ _00257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__09623__A1 _03721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11430__A1 _00514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06615__I _01058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_193_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06988__A2 _01424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11301_ _05801_ _05282_ _05384_ _05393_ _05394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_112_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_154_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_135_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_194_1731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11232_ _01599_ _05140_ _05326_ _05142_ _05327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_84_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11194__B1 _05249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07937__A1 _02161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11163_ as2650.stack\[2\]\[2\] _05212_ _05260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_121_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_36_wb_clk_i clknet_4_6_0_wb_clk_i clknet_leaf_36_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_136_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10114_ _04248_ _04253_ _04266_ _04267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_121_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_1_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06350__I _00798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11094_ _01724_ _05192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_5531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_5553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10045_ as2650.addr_buff\[2\] _04199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_27_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09661__I _03743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07165__A2 _00558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_91_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_79_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11249__A1 _05340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07181__I _01618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11996_ _00365_ clknet_leaf_19_wb_clk_i as2650.r0\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_17_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08114__A1 as2650.stack\[0\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10947_ _05045_ _05047_ _05048_ _04904_ _05049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_44_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08665__A2 _02335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10472__A2 _03873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10878_ _04222_ _04949_ _04982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_176_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_157_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09614__A1 _03777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_185_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10224__A2 _04309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11421__A1 _03565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09090__A2 _01212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06979__A2 _00830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_152_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06971_ _01077_ _01409_ _01410_ _01411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_171_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08710_ as2650.stack\[15\]\[1\] _02978_ _02979_ _02980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05922_ _05775_ _05776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09690_ _02848_ _01286_ _03851_ _03852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_66_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07156__A2 _01593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05853_ _05706_ _05707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08641_ _02784_ _02913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_94_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10160__A1 _02552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06903__A2 _01333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08572_ _02844_ _02845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_130_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08105__A1 as2650.stack\[0\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07523_ _01459_ _01954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09853__A1 _03975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08656__A2 _02849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10999__B1 _05097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07454_ _01852_ _01720_ _01887_ _00024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__10463__A2 _04575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06405_ _00476_ _00843_ _00851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_50_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07385_ as2650.stack\[5\]\[9\] _01816_ _01819_ as2650.stack\[4\]\[9\] _01820_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_22_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08408__A2 _02690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11007__A4 _05105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09124_ _03305_ _03334_ _03345_ _03346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_109_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06336_ _00785_ _00786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__11412__A1 as2650.stack\[9\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05890__A2 _05727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06435__I _00880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09081__A2 _01204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07092__A1 as2650.r123\[1\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09055_ _03174_ _03244_ _03278_ _03281_ _03282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_148_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06267_ _00721_ _00722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_191_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_163_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08006_ as2650.stack\[14\]\[3\] _02362_ _02371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_176_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06198_ _05680_ _00652_ _00656_ _00657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XANTENNA__11176__B1 _01937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11928__D _00297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07919__A1 _02302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11176__C2 _01933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_191_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_132_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06198__A3 _00656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06170__I _00628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_8_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09957_ _02126_ _04069_ _04113_ _02606_ _04114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_131_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08908_ _00439_ _03058_ _03152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_131_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11479__A1 _02604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09888_ net62 _01607_ _04046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08839_ _01277_ _03080_ _03084_ _03085_ _03086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_3425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10151__A1 _03721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11850_ _00010_ clknet_leaf_48_wb_clk_i as2650.cycle\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08097__I _02418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10801_ _02621_ _04878_ _04907_ _04554_ _04908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_2757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09844__A1 _04000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11781_ _00164_ clknet_leaf_85_wb_clk_i as2650.stack\[2\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08647__A2 _02909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10454__A2 _00520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10732_ _02557_ _04841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_158_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10663_ _04583_ _04760_ _04762_ _04772_ _04773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_167_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_161_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05881__A2 _05734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10206__A2 _02594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10594_ _02070_ _04597_ _02082_ _04705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09072__A2 _03259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07083__A1 _05781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07083__B2 _05775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09656__I net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08560__I _00594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11215_ as2650.stack\[8\]\[3\] _05226_ _05310_ as2650.stack\[11\]\[3\] _05311_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_123_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput50 net50 la_data_out[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_150_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput61 net61 la_data_out[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput72 net72 la_data_out[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_68_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11146_ _05135_ _05243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10390__A1 _02835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_95_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11077_ _05173_ _05175_ _05176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_5350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10028_ _04181_ _04182_ _04183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_48_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10142__A1 _00810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08886__A2 _03129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_51_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08638__A2 _02908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11979_ _00348_ clknet_leaf_74_wb_clk_i net60 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_166_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06649__A1 _01090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_32_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06255__I _00640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07170_ _01607_ _01608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_145_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06121_ _00579_ _00580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_195_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_173_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10933__C _04606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06052_ _00510_ _00511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_195_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11158__B1 _03782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11110__B _00824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_193_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09811_ _00822_ _03956_ _03970_ _03971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_140_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10381__A1 _03273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09742_ _03886_ _03902_ _03903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_80_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06954_ _01393_ _00962_ _01394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07129__A2 _01486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08326__A1 _02505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05905_ _05758_ _05759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09673_ _03721_ _03834_ _03835_ _03786_ _00295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_67_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08877__A2 _03122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06885_ _00437_ _00656_ _01325_ _01326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_132_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06888__A1 _05727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10240__I _04385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08624_ _02347_ _00769_ _02868_ _02352_ _02896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_54_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05836_ _05686_ _05689_ _05690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_43_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_184_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08555_ net94 _02826_ _02723_ _02828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_78_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09826__A1 _03978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07506_ _01827_ _01937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10436__A2 _01789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08486_ _00784_ _02759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_50_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07437_ as2650.stack\[9\]\[10\] _01869_ _01758_ as2650.stack\[8\]\[10\] as2650.stack\[10\]\[10\]
+ _01870_ _01871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_51_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_4_13_0_wb_clk_i clknet_3_6_0_wb_clk_i clknet_4_13_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_149_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07852__A3 _02249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05863__A2 _05705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07368_ _01100_ _01803_ _01804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_136_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09107_ _03327_ _03329_ _03330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_136_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06319_ _00647_ _00646_ _00770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_109_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07299_ _01734_ _01735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08801__A2 _03041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06812__A1 _01252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_163_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09038_ _01263_ _03267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08380__I _02665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_191_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_163_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11916__CLK clknet_leaf_94_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_190_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_1892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_151_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11020__B _02349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08565__A1 _02834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11000_ _01091_ _02723_ _00679_ _05099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_104_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10372__A1 _03261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06040__A2 _00498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10911__A3 _05013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output51_I net51 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07724__I _01993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10124__A1 _03769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10124__B2 _04275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06879__A1 _01269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11902_ _00271_ clknet_leaf_73_wb_clk_i as2650.stack\[6\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07540__A2 _01832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11833_ _00216_ clknet_leaf_27_wb_clk_i as2650.r123_2\[1\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11624__A1 _03972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10427__A2 _01789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11764_ _00147_ clknet_leaf_94_wb_clk_i as2650.stack\[5\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10715_ as2650.stack\[6\]\[5\] _04542_ _01789_ as2650.stack\[5\]\[5\] _04824_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_92_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11695_ _00078_ clknet_leaf_120_wb_clk_i as2650.stack\[11\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_186_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06075__I _00533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10646_ _04454_ _04747_ _04756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_195_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_155_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_51_wb_clk_i clknet_4_13_0_wb_clk_i clknet_leaf_51_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_10577_ as2650.stack\[9\]\[2\] _01790_ _01794_ as2650.stack\[8\]\[2\] _04689_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__09386__I _03576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10753__C _04418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_182_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08290__I _02547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06803__I _01233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10325__I _04376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08556__A1 _02342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10363__A1 _01139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06031__A2 _00489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11129_ as2650.stack\[10\]\[1\] _05225_ _05226_ as2650.stack\[8\]\[1\] _05174_ _05227_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__11584__C _04062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08308__A1 _02614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10115__A1 _02218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07516__C1 as2650.stack\[11\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11312__B1 _01961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06670_ _00998_ _01114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__09520__A3 _02737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10666__A2 _04774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_188_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08340_ _02525_ _02639_ _02640_ _02642_ _00155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__11615__A1 _02077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10418__A2 _03757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_189_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08271_ _00483_ _01024_ _02580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_33_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07295__A1 net70 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07222_ as2650.r123\[1\]\[7\] _01197_ _01658_ _01207_ _01659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_20_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07153_ _01461_ _01590_ _01591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_118_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06104_ _00525_ _00562_ _00563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_106_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08414__B _02694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07598__A2 _02025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08795__A1 _02376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07084_ _01521_ _01511_ _01522_ _01377_ _01523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_133_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06035_ _00492_ _00493_ _00494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_195_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_160_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08547__A1 _01597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10354__A1 _00715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06022__A2 _00447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07986_ net4 _02340_ _02354_ _00938_ _02355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__07770__A2 _02163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09725_ net33 _03886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_74_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06937_ _05752_ _01218_ _01377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10106__A1 _02218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11303__B1 _05303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11066__I _05164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09656_ net31 _03819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_27_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06868_ _01308_ _01309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xwrapped_as2650_102 io_oeb[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_3_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xwrapped_as2650_113 io_oeb[32] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_08607_ _02874_ _01668_ _02880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_103_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_124 io_out[37] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_167_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05819_ _05672_ _05673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09587_ _03750_ _02747_ _03751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_27_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_135 la_data_out[52] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_70_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xwrapped_as2650_146 io_oeb[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
X_06799_ _01238_ _01239_ _01240_ _01241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_128_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05999__I _00457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_157 la_data_out[42] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XTAP_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08538_ _02810_ _02811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10409__A2 _00705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11606__A1 _05638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11015__B _02806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11082__A2 _05180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_180_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08469_ _00883_ _00832_ _00855_ _02741_ _02742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_141_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10500_ _04611_ _04612_ _04613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_162_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09027__A2 _03257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11480_ _05539_ _05540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_155_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07038__A1 _00996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10431_ _02779_ _04539_ _04544_ _04545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_137_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08786__A1 as2650.stack\[8\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06623__I _00653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09983__B1 _04051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10362_ _04482_ _04484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_139_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10593__A1 _03914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08250__A3 _02556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_191_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06261__A2 _00625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10293_ _01136_ _04428_ _04429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_5_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12032_ _00401_ clknet_leaf_56_wb_clk_i as2650.r123\[3\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_151_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_191_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07210__A1 _05750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06013__A2 _00471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07761__A2 _02163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10648__A2 _04587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_160_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07403__B _01788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11816_ _00199_ clknet_leaf_111_wb_clk_i as2650.stack\[1\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07277__A1 _00785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11747_ _00130_ clknet_leaf_83_wb_clk_i as2650.stack\[7\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10820__A2 _04102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09018__A2 _03101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11678_ _00061_ clknet_leaf_130_wb_clk_i as2650.stack\[12\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07029__A1 _01463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_30_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10629_ _04735_ _04736_ _04739_ _04740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_102_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07629__I _02055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_183_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10055__I net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_142_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08529__A1 _01787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11595__B _04435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_151_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07201__A1 _05742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07840_ _02239_ _02207_ _02243_ _02241_ _00054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_69_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09741__A3 net93 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07752__A2 _02149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07771_ _02128_ _02184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_56_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09510_ _00622_ _00911_ _03640_ _03675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_42_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06722_ _01090_ _00592_ _01092_ _01165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_80_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07504__A2 _01933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_40_wb_clk_i_I clknet_4_6_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09441_ as2650.stack\[5\]\[0\] _03615_ _03616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06653_ _01076_ _01079_ _01095_ _01072_ _01096_ _01097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
XFILLER_25_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08195__I _02213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09372_ as2650.stack\[3\]\[5\] _03552_ _03566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06584_ net50 _01028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__11761__CLK clknet_leaf_82_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08323_ _02138_ _02630_ _02631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_32_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08254_ _02562_ _00850_ _02550_ _02563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_21_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07205_ _01547_ _01551_ _01642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06491__A2 _00872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08185_ _02507_ _02508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_174_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08768__A1 _02151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08144__B _02474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07136_ _01572_ _01567_ _01574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10575__A1 _02789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07067_ _01375_ _01382_ _01506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06243__A2 _00699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06018_ _05684_ _00477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07991__A2 _02000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10327__A1 _00736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10878__A2 _04949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07743__A2 _02161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07969_ _02334_ _02337_ _02338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09708_ _00638_ _03870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10980_ _05079_ _05080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_28_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09496__A2 _00694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09639_ _03797_ _03763_ _03801_ _03802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_28_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_164_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09248__A2 _03465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11601_ _05608_ _05644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_93_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_93_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11532_ _01986_ _05177_ _05580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__08833__I _03079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10802__A2 _04906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_183_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06482__A2 _00925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11463_ _01022_ _05672_ _05522_ _05523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_139_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07449__I _01777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08759__A1 as2650.stack\[1\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10414_ _04323_ _04520_ _04523_ _04527_ _04528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_165_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10566__A1 _04668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11394_ as2650.stack\[9\]\[14\] _05456_ _05471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_136_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10345_ _04468_ _00334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_87_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_139_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10276_ _04400_ _00822_ _04412_ _04414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_105_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10318__A1 _03609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11634__CLK clknet_leaf_37_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12015_ _00384_ clknet_leaf_100_wb_clk_i as2650.stack\[9\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10869__A2 _04789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06537__A3 _00980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_171_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09487__A2 _02348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11784__CLK clknet_leaf_85_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07498__A1 _01449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11294__A2 _05386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_124_wb_clk_i_I clknet_4_0_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08743__I _02693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08462__A3 _00982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06473__A2 _00811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10006__B1 _04160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07359__I _01794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06263__I _00714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10557__A1 net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09411__A2 _03589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_7_wb_clk_i_I clknet_4_4_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10021__A3 _04126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09990_ _04142_ _04144_ _04145_ _04146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_89_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10941__C _03816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_130_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08941_ _01460_ _03112_ _03182_ _03087_ _03183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_131_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05984__A1 _05703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09175__A1 _05758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10513__I _04540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08872_ _01150_ _03113_ _03117_ _03085_ _03118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_111_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07823_ _01518_ _02190_ _02124_ _02229_ _02230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_57_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07754_ _02170_ _02156_ _02164_ _02171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_56_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10669__B _01775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07822__I net69 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06705_ _01146_ _01147_ _01148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_53_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11285__A2 _05370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07685_ _01954_ _02084_ _02108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_148_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08150__A2 _02480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09424_ as2650.ivec\[2\] _03267_ _03604_ _03605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06438__I _00663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06636_ _00663_ _01080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_13_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06161__A1 _00529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09355_ _02651_ _03553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11037__A2 _04553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06567_ _01010_ _01011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_100_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08306_ _02341_ _02336_ _02615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_51_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08989__A1 _03028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11588__A3 _02965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09286_ _02670_ _03500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_165_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06498_ _00940_ _00941_ _00942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__10796__A1 _03820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08237_ _00898_ _00615_ _02546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_14_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07661__A1 _02082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_181_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_153_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06173__I _00631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08168_ _02318_ _02489_ _02494_ _02496_ _00129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_140_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10548__A1 _03876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_194_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_108_wb_clk_i clknet_4_3_0_wb_clk_i clknet_leaf_108_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_146_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11657__CLK clknet_leaf_124_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07119_ _01556_ _01557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__07413__A1 _01203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06216__A2 _00644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08099_ _02384_ _02436_ _02441_ _02443_ _00113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_49_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10130_ _04250_ _04230_ _04281_ _04282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_161_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06901__I _01331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_192_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10061_ _04142_ _04169_ _04215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_5724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_134_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06519__A3 _00962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07716__A2 _01993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08828__I _03057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10963_ _05025_ _05040_ _05064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__11276__A2 _05366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10323__I1 as2650.holding_reg\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08141__A2 _02468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10894_ as2650.ivec\[5\] _04972_ _04941_ _04975_ _04873_ _04998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_43_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11028__A2 _01019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11579__A3 _02965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08563__I _01565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09641__A2 _03092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10787__A1 _04879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_180_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11515_ _02856_ _02770_ _05563_ _05564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_157_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06455__A2 _00557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11446_ _01889_ _05499_ _05504_ as2650.r123\[2\]\[3\] _05511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_171_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_158_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11377_ _05459_ _05460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_140_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07955__A2 _02279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10328_ _04456_ _04457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10259_ _04401_ _00315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05981__A4 _00439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10711__A1 _03642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08738__I _02688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07470_ _01897_ _01898_ _01902_ _01903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__06143__A1 _00601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06421_ _00866_ _00763_ _00849_ _00867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__07891__A1 _02276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_124_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09140_ _05759_ _01516_ _03362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_148_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06352_ _00800_ _00801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_147_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09071_ _03214_ _03257_ _03294_ _03295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_147_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06283_ _00736_ _00737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_30_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08022_ as2650.stack\[14\]\[7\] _02360_ _02356_ _02383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_129_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08422__B _02701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09973_ _03948_ _04129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_89_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10950__A1 _01926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10950__B2 _03666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08924_ _03165_ _03151_ _03080_ _03166_ _03167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_150_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09699__A2 _01271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08855_ _00835_ _03101_ _03102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_4319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07806_ _02189_ _02214_ _02215_ _02210_ _00048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__08371__A2 _02649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08786_ as2650.stack\[8\]\[3\] _03026_ _03038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05998_ _05720_ _00454_ _00456_ _00457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_85_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07737_ _02139_ _02157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_72_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11258__A2 _00873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08123__A2 _02425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06168__I _00626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06134__A1 _00590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07668_ _02046_ _02092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_81_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09407_ as2650.stack\[6\]\[5\] _03585_ _03574_ _03593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06619_ _05720_ _05777_ _05778_ _05708_ _01063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_13_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06685__A2 _00979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07882__A1 _02272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07599_ _01771_ _02027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09479__I _00541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08383__I _02213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09338_ _03239_ _02634_ _03518_ _03539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_90_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10769__A1 _02115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_178_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11023__B _02742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07634__A1 _02053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09269_ _03475_ _03484_ _03485_ _00241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11430__A2 _00997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11300_ _02837_ _05205_ _05392_ _05393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_153_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_159_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09387__A1 as2650.stack\[6\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11231_ _01431_ _05138_ _05325_ _02960_ _05326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_107_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11194__A1 _03148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08332__B _02633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07727__I _02022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07937__A2 _02237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11162_ _05209_ _05256_ _05258_ _05259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_134_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10113_ _02218_ _04111_ _04265_ _03830_ _04266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_96_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11093_ net79 _02589_ _05191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_5521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09942__I _03733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10044_ _04068_ _04197_ _04198_ _00303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_76_wb_clk_i clknet_4_11_0_wb_clk_i clknet_leaf_76_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_5576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11995_ _00364_ clknet_leaf_26_wb_clk_i as2650.r0\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_16_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08114__A2 _02440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_182_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_188_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06125__A1 _00556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10946_ _04226_ _05028_ _05048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_90_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07873__A1 as2650.stack\[12\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10877_ _04808_ _04978_ _04980_ _04891_ _04981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_176_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_31_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09614__A2 _03731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10328__I _04456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11421__A2 _05487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_195_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_1518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11972__CLK clknet_leaf_39_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09378__A1 _03568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11429_ _05496_ _03337_ _05497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_126_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11587__C _05076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06541__I as2650.cycle\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10932__A1 _04604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06600__A2 _00946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06970_ _01406_ _01408_ _01397_ _01410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_113_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input5_I io_in[33] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05921_ _05774_ _05775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_140_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09550__A1 _02552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08640_ _02907_ _02910_ _02911_ _02912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_05852_ as2650.ins_reg\[1\] _05705_ _05706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__07372__I as2650.r123\[0\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10160__A2 _00555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08571_ _01043_ _02844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_82_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_35_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08105__A2 _02440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09302__A1 _02376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07522_ _01939_ _01946_ _01952_ _01883_ _01953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_58_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10999__A1 _02841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09853__A2 _02955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10999__B2 _00951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_180_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07453_ _01295_ _01722_ _01853_ _01886_ _01887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__10463__A3 _04576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06404_ _00514_ _00849_ _00845_ _00850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_07384_ _01818_ _01819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09123_ _03308_ _03333_ _03345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_148_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06335_ _00784_ _00785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07616__A1 _02039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11412__A2 _05478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09081__A3 _01637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09054_ _03279_ _03262_ _03280_ _03281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_135_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_178_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06266_ _00531_ as2650.cycle\[10\] _00721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_190_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_175_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_194_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08005_ _02067_ _02357_ _02369_ _02370_ _00092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__09369__A1 _02456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06197_ _00655_ _00656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_11_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11176__A1 as2650.stack\[8\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08152__B _02481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_191_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07919__A2 _02297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11176__B2 as2650.stack\[11\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_172_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09956_ _04091_ _04095_ _04112_ _04113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_63_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08907_ _03058_ _03151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_4105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09887_ _00718_ _04040_ _04044_ _04004_ _04045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_4116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11479__A2 _05537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09541__A1 _00891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08838_ _03077_ _03085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06355__A1 _00671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11018__B _03745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08769_ _02022_ _03024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11845__CLK clknet_leaf_54_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10800_ _02571_ _02924_ _04907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06107__A1 _00563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11780_ _00163_ clknet_leaf_93_wb_clk_i as2650.stack\[3\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11100__A1 _03148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10857__B _04186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10731_ _04790_ _04793_ _04839_ _00732_ _04840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_92_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07855__A1 as2650.stack\[12\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10454__A3 _00894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10662_ _04609_ _04748_ _04770_ _04771_ _04772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__11995__CLK clknet_leaf_26_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_185_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_123_wb_clk_i clknet_4_2_0_wb_clk_i clknet_leaf_123_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_103_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07607__A1 _02030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10593_ _03914_ _04653_ _04704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_194_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10757__A4 _04864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06361__I _00627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11214_ _01879_ _05310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_141_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput40 net40 io_out[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__10914__A1 _04242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput51 net51 la_data_out[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_155_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09780__A1 _02858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput62 net62 la_data_out[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_11145_ _02814_ _00842_ _05242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xoutput73 net73 la_data_out[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_110_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06594__A1 _00489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11076_ as2650.stack\[10\]\[0\] _01959_ _01936_ as2650.stack\[8\]\[0\] _05174_ _05175_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XTAP_5351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09532__A1 _05697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10027_ net38 _04133_ _04182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_3_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10142__A2 _04293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06897__A2 _01239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08099__A1 _02384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11978_ _00347_ clknet_leaf_74_wb_clk_i net58 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_147_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09835__A2 _03993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06649__A2 _00592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10929_ _02224_ _02216_ _05000_ _05031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__07846__A1 _02053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_71_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12000__CLK clknet_4_10_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_53_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_34_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06120_ _00578_ _00559_ _00579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_121_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08271__A1 _00483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11598__B _05635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_172_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06051_ _05676_ _00510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_133_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11158__A1 _00426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11158__B2 _05240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11718__CLK clknet_leaf_134_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08023__A1 _02122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10905__A1 _02212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09810_ _02094_ _03725_ _03916_ _03969_ _03883_ _03970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_113_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09771__A1 _00728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09582__I _03745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09741_ net32 net31 net93 _03902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_101_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06953_ _05760_ _01393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05904_ as2650.r0\[4\] _05758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_95_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09672_ _03819_ _03720_ _03835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_67_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06884_ as2650.holding_reg\[3\] _00829_ _01325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_95_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08623_ _02776_ _02892_ _02895_ _00185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_67_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05835_ _05687_ _05688_ _05689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__06888__A2 _00988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08554_ _02596_ _02827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_54_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07505_ _01830_ _01936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_74_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07837__A1 _02239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08485_ _00798_ _00615_ _02758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_35_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07436_ _01746_ _01870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_74_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_50_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07367_ _01726_ _01803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09106_ _03310_ _03328_ _03329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__08661__I net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06318_ _00768_ _00769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_191_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07298_ _01733_ _01734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_191_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_121_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09037_ _03266_ _00228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11301__B _05384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06812__A2 _01123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06249_ _00700_ _00705_ _00706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_69_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11149__A1 _02135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08014__A1 _02376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08565__A2 _02835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09762__A1 _03734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09706__B _00679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09939_ _04049_ _04055_ _04047_ _04096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_77_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11527__I _05570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output44_I net44 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11901_ _00270_ clknet_leaf_73_wb_clk_i as2650.stack\[6\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_111_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_172_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06879__A2 _01284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11832_ _00215_ clknet_leaf_27_wb_clk_i as2650.r123_2\[1\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12023__CLK clknet_leaf_38_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11763_ _00146_ clknet_leaf_80_wb_clk_i as2650.stack\[5\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10714_ as2650.stack\[7\]\[5\] _04822_ _01793_ as2650.stack\[4\]\[5\] _04823_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06356__I _00601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11694_ _00077_ clknet_leaf_119_wb_clk_i as2650.stack\[11\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_14_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_161_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10645_ _03958_ _02955_ _04754_ _04755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_35_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09667__I _00451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08571__I _01043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08253__A1 _00472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10576_ _02780_ _04684_ _04687_ _04688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_154_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06091__I as2650.cycle\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08005__A1 _02067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_91_wb_clk_i clknet_4_8_0_wb_clk_i clknet_leaf_91_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__08556__A2 _02826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_20_wb_clk_i clknet_4_5_0_wb_clk_i clknet_leaf_20_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_111_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11560__A1 _05599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11128_ _01816_ _05226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_3_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09505__A1 _01091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08308__A2 _02616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_5170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06319__A1 _00647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11059_ _02131_ _01990_ _05158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_5181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10115__A2 _03788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07516__B1 _01941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11312__A1 as2650.stack\[14\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07516__C2 _01940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11312__B2 as2650.stack\[12\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_30_wb_clk_i_I clknet_4_7_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09520__A4 _03672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11076__B1 _01936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11172__I _01900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08270_ _02571_ _02573_ _02576_ _02578_ _02579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__08492__A1 _02764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07221_ _01626_ _01657_ _01658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_32_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11379__A1 _02663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07152_ _05802_ _05807_ _01423_ _01590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__08244__A1 _02552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10051__A1 _04175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06103_ _00531_ _00561_ _00562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_161_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08795__A2 _03029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07083_ _05781_ _01362_ _01380_ _05775_ _01522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_172_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06034_ _05788_ _00493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_82_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08547__A2 _01459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09744__A1 _00633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10354__A2 _00906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11551__A1 _03657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07985_ _02338_ _02344_ _02353_ _00853_ _02354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_59_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09724_ _00728_ _03885_ _00296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06936_ _01357_ _01362_ _01376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_151_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10106__A2 _04101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07507__B1 _01937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11303__A1 as2650.stack\[5\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11303__B2 as2650.stack\[7\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09655_ _03816_ _03817_ _03818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_28_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06867_ _05807_ _01308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_55_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05908__I1 as2650.r123\[0\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xwrapped_as2650_103 io_oeb[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_08606_ _01581_ _02877_ _02878_ _01416_ _02879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_43_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xwrapped_as2650_114 io_out[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_55_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05818_ _05671_ _05672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09586_ _00778_ _03750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_125 la_data_out[33] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__06730__A1 _01171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06798_ _01238_ _01239_ _00839_ _01240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_136 la_data_out[54] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xwrapped_as2650_147 io_oeb[33] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
X_08537_ _02764_ _02810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_158 la_data_out[44] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XANTENNA__11067__B1 _01942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10409__A3 _04521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11606__A2 _04443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_169_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10200__B _00525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08468_ _05671_ _02740_ _02741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__08483__A1 _02754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_195_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07419_ _01718_ _01853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08399_ as2650.stack\[2\]\[14\] _02666_ _02687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_195_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10854__C _04891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10430_ _04540_ _04541_ _04543_ _04544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_195_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07038__A2 _01458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08235__A1 as2650.stack\[5\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10042__A1 _02205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09983__A1 _02125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08786__A2 _03026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10361_ _04482_ _04483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_163_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06125__B _00572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10593__A2 _04653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08250__A4 _02558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06261__A3 _00715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10292_ _02349_ _04428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_105_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12031_ _00400_ clknet_leaf_59_wb_clk_i as2650.r123\[3\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_156_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06549__A1 _00992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08340__B _02640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11542__A1 _01773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07210__A2 _01515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08710__A2 _02978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06721__A1 _00996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_146_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11815_ _00198_ clknet_leaf_111_wb_clk_i as2650.stack\[1\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_114_wb_clk_i_I clknet_4_2_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07277__A2 _00974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11746_ _00129_ clknet_leaf_113_wb_clk_i as2650.stack\[7\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_186_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11677_ _00060_ clknet_leaf_130_wb_clk_i as2650.stack\[12\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_15_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10764__C _00732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08226__A1 _02516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10628_ _01733_ _04737_ _04738_ _04739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_174_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10033__A1 _03824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09974__A1 _04024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10336__I _00750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_182_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10559_ _03790_ _05782_ _04671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_154_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09974__B2 _04129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06788__A1 _01227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07985__B1 _02353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10584__A2 _04695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10780__B _04608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07645__I _02070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11533__A1 _01262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07201__A2 _01198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11167__I _00755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10071__I _00982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07770_ as2650.stack\[11\]\[7\] _02163_ _02183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_37_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06721_ _00996_ _01127_ _01163_ _01164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_133_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09440_ _03614_ _03615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06652_ _01093_ _01096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_1724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07380__I _01814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09371_ _02100_ _03565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06583_ _01025_ _01026_ _01027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_1779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08322_ _01934_ _01769_ _02630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_178_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08465__A1 _02582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08253_ _00472_ _00834_ _02562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10447__S _00441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07204_ _01639_ _01640_ _01641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__08217__A1 _01985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06724__I _00664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08184_ _02506_ _02507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10246__I _04384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09965__A1 _04118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07135_ _01572_ _01567_ _01573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__08768__A2 _02480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11221__B1 _05306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07066_ _01383_ _01384_ _01505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10690__B _04570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06017_ _05688_ _00476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__09717__A1 _03752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07991__A3 _02272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10327__A2 _04455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07555__I _01030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07968_ _02336_ _02337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_74_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06951__A1 _01390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06919_ _01359_ _01360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09707_ _00630_ _03865_ _03868_ _03728_ _03869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_07899_ as2650.stack\[10\]\[2\] _02274_ _02288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_74_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09638_ _03762_ _03800_ _03801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_112_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09569_ _00793_ _03733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_31_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11600_ _05643_ _00414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_58_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08456__A1 _02725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_180_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10865__B _04969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11531_ _02777_ _05579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10263__A1 _00568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_36_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10802__A3 _04908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_141_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08208__A1 as2650.stack\[6\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11462_ _00859_ _05522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_137_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09956__A1 _04091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10413_ _04524_ _04525_ _04308_ _04526_ _04527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__08759__A2 _03004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11212__B1 _05269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_183_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_164_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11393_ _02684_ _05467_ _05468_ _05470_ _00380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_136_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09945__I _00688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10566__A2 _04648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10344_ _00811_ _00751_ _04458_ _00825_ _04468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_87_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10275_ _01121_ _04412_ _04413_ _04405_ _00319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_155_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10318__A2 _02903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11515__A1 _02856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12014_ _00383_ clknet_leaf_90_wb_clk_i as2650.stack\[9\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_78_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07195__A1 _01541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11929__CLK clknet_leaf_62_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06809__I _01250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09892__B1 _01464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05902__C1 _05755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07133__C _00666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10775__B _04802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10254__A1 _00978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11729_ _00112_ clknet_leaf_88_wb_clk_i as2650.stack\[0\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10494__C _04606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10006__A1 _04135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10006__B2 _04161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11203__B1 _05297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10557__A2 _05754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_131_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_170_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08940_ _03179_ _03181_ _03085_ _03182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_143_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10309__A2 _04441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11506__A1 _04948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05984__A2 _00442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07375__I _01809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09175__A2 _02233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08871_ _01146_ _03114_ _03116_ _03117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_48_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07822_ net69 _02229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_57_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06933__A1 _05766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_69_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07753_ _02086_ _02170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_42_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06704_ _00932_ _01147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_38_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07684_ _02106_ _02107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07489__A2 _01865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09423_ _03600_ _03604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_06635_ _01077_ _01078_ _01079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_168_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09354_ _03545_ _03552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06566_ _01008_ _01009_ _01010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__08438__A1 _02675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06882__C _01250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08305_ _02613_ _02614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09285_ _02976_ _02681_ _03499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07110__A1 _05750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06497_ _00478_ _00941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_138_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10796__A2 _00689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08236_ _02527_ _02541_ _02542_ _02545_ _00148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_53_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06464__A3 _00580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09938__A1 _00717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08167_ as2650.stack\[7\]\[9\] _02495_ _02496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_146_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10548__A2 _03866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07118_ _05732_ _01199_ _01556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08098_ _02276_ _02442_ _02431_ _02443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_106_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07049_ _01487_ _01488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_106_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07285__I _01099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09166__A2 _03363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10060_ _04170_ _04213_ _04214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_5714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06924__A1 _01361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_169_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08677__A1 _02938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10962_ _01155_ _05062_ _02331_ _05063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_95_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10484__A1 net90 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10893_ _03662_ _04975_ _04994_ _04996_ _03832_ _04997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_44_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_77_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08429__A1 _02133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11270__I _05159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_157_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11514_ _05561_ _05558_ _05562_ _05563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__06364__I _00810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11203__C _05298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11445_ _05496_ _03431_ _05510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_172_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_165_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09675__I _03719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11376_ _02465_ _02138_ _05459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_124_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10327_ _00736_ _04455_ _00507_ _04456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_152_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11751__CLK clknet_leaf_88_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10258_ _04399_ _04400_ _04385_ _04401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_112_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07168__A1 _05801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10189_ _00560_ _00565_ _04338_ _04339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_117_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10711__A2 _04810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07923__I _02157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_187_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_47_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06143__A2 _05702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06420_ _00651_ _00866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_34_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07891__A2 _02279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06351_ _00799_ _00800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09070_ _01980_ _03251_ _03278_ _03294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_148_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06274__I _00727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06282_ _00735_ _00736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_120_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08021_ _02381_ _02365_ _02382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09585__I _02865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10952__C _04643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_fanout93_I net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09972_ _04116_ _04127_ _04128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_170_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10950__A2 _04622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08923_ _05813_ _03151_ _03166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_103_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08854_ _01103_ _03100_ _03101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06906__A1 _01081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07805_ as2650.stack\[14\]\[10\] _02208_ _02215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08371__A3 _02664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08785_ _02077_ _03037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05997_ _00455_ _05679_ _00456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_73_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11355__I _05446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07736_ _02155_ _02156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_38_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06449__I _00894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10466__A1 _03726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07667_ _02090_ _02091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_129_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06134__A2 _00592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07331__A1 as2650.stack\[2\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06618_ _01015_ _00665_ _01062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09406_ _02177_ _03579_ _03592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07598_ as2650.stack\[13\]\[0\] _02025_ _02026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07882__A2 _02146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10218__A1 _00789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06549_ _00992_ _00544_ _00993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_51_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09337_ as2650.stack\[4\]\[6\] _03526_ _03538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10769__A2 _04007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09268_ _03202_ _03338_ _03340_ as2650.r123_2\[2\]\[6\] _03485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_142_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07634__A2 _02060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08219_ _02534_ _02535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_177_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09199_ _05731_ _02233_ _03419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_147_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09495__I _03661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11230_ _05129_ _02223_ _05324_ _02818_ _05325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__11774__CLK clknet_leaf_82_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09387__A2 _03577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07398__A1 as2650.stack\[3\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11194__A2 _02815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_150_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11161_ as2650.stack\[5\]\[2\] _05257_ _05223_ as2650.stack\[7\]\[2\] as2650.stack\[6\]\[2\]
+ _02387_ _05258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_162_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output74_I net74 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10112_ _04109_ _04259_ _04263_ _04264_ _04265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__10941__A2 _05028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11092_ _00805_ _00431_ _05190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_5511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10043_ _04181_ _03976_ _04165_ _04198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_5544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_5555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06373__A2 _00816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_99_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11994_ _00363_ clknet_4_5_0_wb_clk_i as2650.r0\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_99_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10457__A1 _05777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10945_ _04897_ _05046_ _05047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_95_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08574__I _02846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10876_ _04708_ _04979_ _04980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07873__A2 _02260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10209__A1 _03684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_188_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_164_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09619__B _03780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07918__I _02128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09378__A2 _03562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11428_ _01107_ _05496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06822__I _01051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11359_ _05448_ _00368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_153_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_152_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10932__A2 _05033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06600__A3 _00927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05920_ as2650.r0\[0\] _05774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_67_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07653__I _02077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05851_ as2650.ins_reg\[0\] _05705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_13_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08570_ _00630_ _02842_ _02843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_66_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07521_ _01947_ _01948_ _01951_ _01952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09302__A2 _03502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_184_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06116__A2 _00561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08510__B1 _01780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10947__C _04904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10999__A2 _02772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07452_ _01728_ _01884_ _01885_ _01849_ _01886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_161_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05875__A1 _05724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06403_ _00667_ _00849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_182_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09066__A1 _01974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07383_ _01817_ _01818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_91_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09122_ _03300_ _03336_ _03343_ _03344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_124_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06334_ _00559_ _00784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08813__A1 _00953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11797__CLK clknet_leaf_120_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09053_ _01926_ _03250_ _03280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_124_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10620__A1 _01734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06265_ as2650.cycle\[2\] _00720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_175_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09529__B _02549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07828__I _02233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08004_ as2650.stack\[14\]\[2\] _02360_ _02366_ _02370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_159_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06196_ _00654_ _00655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_117_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11176__A2 _01914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_171_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09955_ _03830_ _04110_ _04111_ _02126_ _04112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_106_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08906_ _01310_ _03150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_4106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08659__I net77 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09886_ _03811_ _04043_ _04044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09541__A2 _02005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08837_ _00428_ _03082_ _03079_ _03083_ _03084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_3405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07552__A1 _01980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06179__I _00637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11018__C _00647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08768_ _02151_ _02480_ _03023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_26_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10439__A1 _04545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07719_ _02133_ _02137_ _02138_ _02139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_57_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06107__A2 _00565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_4_0_0_wb_clk_i_I clknet_3_0_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11960__D _00329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08699_ _02969_ _02970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11100__A2 _02833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10730_ _04821_ _04838_ _04839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_92_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_158_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10661_ _04332_ _04771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11034__B _02724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_107_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10592_ _03914_ _04646_ _04703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__08804__A1 as2650.stack\[8\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10206__A4 _04355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10611__A1 _03960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07738__I _02157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06642__I _00593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_182_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11213_ _05307_ _05308_ _05309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_135_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput30 net30 io_out[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput41 net41 io_out[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_162_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10914__A2 _04987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput52 net52 la_data_out[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_68_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11144_ _00594_ _05241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09780__A2 _01429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput63 net63 la_data_out[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_96_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xoutput74 net74 la_data_out[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__06798__B _00839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06594__A2 _01037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07791__A1 as2650.stack\[14\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_172_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11075_ _05164_ _05174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_163_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10127__B1 _04278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08569__I _02841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10026_ net39 _04181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_114_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10678__A1 _04532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_188_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09532__A2 _00840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06346__A2 _00586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_20_wb_clk_i_I clknet_4_5_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06346__B3 _00795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06089__I _00536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08099__A2 _02436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09296__A1 _03037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11977_ _00346_ clknet_leaf_74_wb_clk_i net57 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_17_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10767__C _00739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06649__A3 _01092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10928_ _05026_ _04228_ _05029_ _05030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07846__A2 _02227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09048__A1 _03162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10859_ _04794_ _04961_ _04962_ _04963_ _04964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_13_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10602__A1 _04709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08271__A2 _01024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07648__I _02073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06050_ _00502_ _00508_ _00509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_172_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_172_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11158__A2 _00680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08023__A2 _02373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10905__A2 _04949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09740_ _03893_ _03900_ _03793_ _03901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_141_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06952_ as2650.holding_reg\[4\] _00665_ _01391_ _01392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_119_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
.ends

