magic
tech gf180mcuD
magscale 1 5
timestamp 1700058980
<< obsm1 >>
rect 672 1538 79296 58438
<< metal2 >>
rect 2576 59600 2632 60000
rect 4592 59600 4648 60000
rect 6608 59600 6664 60000
rect 8624 59600 8680 60000
rect 10640 59600 10696 60000
rect 12656 59600 12712 60000
rect 14672 59600 14728 60000
rect 16688 59600 16744 60000
rect 18704 59600 18760 60000
rect 20720 59600 20776 60000
rect 22736 59600 22792 60000
rect 24752 59600 24808 60000
rect 26768 59600 26824 60000
rect 28784 59600 28840 60000
rect 30800 59600 30856 60000
rect 32816 59600 32872 60000
rect 34832 59600 34888 60000
rect 36848 59600 36904 60000
rect 38864 59600 38920 60000
rect 40880 59600 40936 60000
rect 42896 59600 42952 60000
rect 44912 59600 44968 60000
rect 46928 59600 46984 60000
rect 48944 59600 49000 60000
rect 50960 59600 51016 60000
rect 52976 59600 53032 60000
rect 54992 59600 55048 60000
rect 57008 59600 57064 60000
rect 59024 59600 59080 60000
rect 61040 59600 61096 60000
rect 63056 59600 63112 60000
rect 65072 59600 65128 60000
rect 67088 59600 67144 60000
rect 69104 59600 69160 60000
rect 71120 59600 71176 60000
rect 73136 59600 73192 60000
rect 75152 59600 75208 60000
rect 77168 59600 77224 60000
rect 336 0 392 400
rect 1120 0 1176 400
rect 1904 0 1960 400
rect 2688 0 2744 400
rect 3472 0 3528 400
rect 4256 0 4312 400
rect 5040 0 5096 400
rect 5824 0 5880 400
rect 6608 0 6664 400
rect 7392 0 7448 400
rect 8176 0 8232 400
rect 8960 0 9016 400
rect 9744 0 9800 400
rect 10528 0 10584 400
rect 11312 0 11368 400
rect 12096 0 12152 400
rect 12880 0 12936 400
rect 13664 0 13720 400
rect 14448 0 14504 400
rect 15232 0 15288 400
rect 16016 0 16072 400
rect 16800 0 16856 400
rect 17584 0 17640 400
rect 18368 0 18424 400
rect 19152 0 19208 400
rect 19936 0 19992 400
rect 20720 0 20776 400
rect 21504 0 21560 400
rect 22288 0 22344 400
rect 23072 0 23128 400
rect 23856 0 23912 400
rect 24640 0 24696 400
rect 25424 0 25480 400
rect 26208 0 26264 400
rect 26992 0 27048 400
rect 27776 0 27832 400
rect 28560 0 28616 400
rect 29344 0 29400 400
rect 30128 0 30184 400
rect 30912 0 30968 400
rect 31696 0 31752 400
rect 32480 0 32536 400
rect 33264 0 33320 400
rect 34048 0 34104 400
rect 34832 0 34888 400
rect 35616 0 35672 400
rect 36400 0 36456 400
rect 37184 0 37240 400
rect 37968 0 38024 400
rect 38752 0 38808 400
rect 39536 0 39592 400
rect 40320 0 40376 400
rect 41104 0 41160 400
rect 41888 0 41944 400
rect 42672 0 42728 400
rect 43456 0 43512 400
rect 44240 0 44296 400
rect 45024 0 45080 400
rect 45808 0 45864 400
rect 46592 0 46648 400
rect 47376 0 47432 400
rect 48160 0 48216 400
rect 48944 0 49000 400
rect 49728 0 49784 400
rect 50512 0 50568 400
rect 51296 0 51352 400
rect 52080 0 52136 400
rect 52864 0 52920 400
rect 53648 0 53704 400
rect 54432 0 54488 400
rect 55216 0 55272 400
rect 56000 0 56056 400
rect 56784 0 56840 400
rect 57568 0 57624 400
rect 58352 0 58408 400
rect 59136 0 59192 400
rect 59920 0 59976 400
rect 60704 0 60760 400
rect 61488 0 61544 400
rect 62272 0 62328 400
rect 63056 0 63112 400
rect 63840 0 63896 400
rect 64624 0 64680 400
rect 65408 0 65464 400
rect 66192 0 66248 400
rect 66976 0 67032 400
rect 67760 0 67816 400
rect 68544 0 68600 400
rect 69328 0 69384 400
rect 70112 0 70168 400
rect 70896 0 70952 400
rect 71680 0 71736 400
rect 72464 0 72520 400
rect 73248 0 73304 400
rect 74032 0 74088 400
rect 74816 0 74872 400
rect 75600 0 75656 400
rect 76384 0 76440 400
rect 77168 0 77224 400
rect 77952 0 78008 400
rect 78736 0 78792 400
rect 79520 0 79576 400
<< obsm2 >>
rect 350 59570 2546 59600
rect 2662 59570 4562 59600
rect 4678 59570 6578 59600
rect 6694 59570 8594 59600
rect 8710 59570 10610 59600
rect 10726 59570 12626 59600
rect 12742 59570 14642 59600
rect 14758 59570 16658 59600
rect 16774 59570 18674 59600
rect 18790 59570 20690 59600
rect 20806 59570 22706 59600
rect 22822 59570 24722 59600
rect 24838 59570 26738 59600
rect 26854 59570 28754 59600
rect 28870 59570 30770 59600
rect 30886 59570 32786 59600
rect 32902 59570 34802 59600
rect 34918 59570 36818 59600
rect 36934 59570 38834 59600
rect 38950 59570 40850 59600
rect 40966 59570 42866 59600
rect 42982 59570 44882 59600
rect 44998 59570 46898 59600
rect 47014 59570 48914 59600
rect 49030 59570 50930 59600
rect 51046 59570 52946 59600
rect 53062 59570 54962 59600
rect 55078 59570 56978 59600
rect 57094 59570 58994 59600
rect 59110 59570 61010 59600
rect 61126 59570 63026 59600
rect 63142 59570 65042 59600
rect 65158 59570 67058 59600
rect 67174 59570 69074 59600
rect 69190 59570 71090 59600
rect 71206 59570 73106 59600
rect 73222 59570 75122 59600
rect 75238 59570 77138 59600
rect 77254 59570 79562 59600
rect 350 430 79562 59570
rect 422 345 1090 430
rect 1206 345 1874 430
rect 1990 345 2658 430
rect 2774 345 3442 430
rect 3558 345 4226 430
rect 4342 345 5010 430
rect 5126 345 5794 430
rect 5910 345 6578 430
rect 6694 345 7362 430
rect 7478 345 8146 430
rect 8262 345 8930 430
rect 9046 345 9714 430
rect 9830 345 10498 430
rect 10614 345 11282 430
rect 11398 345 12066 430
rect 12182 345 12850 430
rect 12966 345 13634 430
rect 13750 345 14418 430
rect 14534 345 15202 430
rect 15318 345 15986 430
rect 16102 345 16770 430
rect 16886 345 17554 430
rect 17670 345 18338 430
rect 18454 345 19122 430
rect 19238 345 19906 430
rect 20022 345 20690 430
rect 20806 345 21474 430
rect 21590 345 22258 430
rect 22374 345 23042 430
rect 23158 345 23826 430
rect 23942 345 24610 430
rect 24726 345 25394 430
rect 25510 345 26178 430
rect 26294 345 26962 430
rect 27078 345 27746 430
rect 27862 345 28530 430
rect 28646 345 29314 430
rect 29430 345 30098 430
rect 30214 345 30882 430
rect 30998 345 31666 430
rect 31782 345 32450 430
rect 32566 345 33234 430
rect 33350 345 34018 430
rect 34134 345 34802 430
rect 34918 345 35586 430
rect 35702 345 36370 430
rect 36486 345 37154 430
rect 37270 345 37938 430
rect 38054 345 38722 430
rect 38838 345 39506 430
rect 39622 345 40290 430
rect 40406 345 41074 430
rect 41190 345 41858 430
rect 41974 345 42642 430
rect 42758 345 43426 430
rect 43542 345 44210 430
rect 44326 345 44994 430
rect 45110 345 45778 430
rect 45894 345 46562 430
rect 46678 345 47346 430
rect 47462 345 48130 430
rect 48246 345 48914 430
rect 49030 345 49698 430
rect 49814 345 50482 430
rect 50598 345 51266 430
rect 51382 345 52050 430
rect 52166 345 52834 430
rect 52950 345 53618 430
rect 53734 345 54402 430
rect 54518 345 55186 430
rect 55302 345 55970 430
rect 56086 345 56754 430
rect 56870 345 57538 430
rect 57654 345 58322 430
rect 58438 345 59106 430
rect 59222 345 59890 430
rect 60006 345 60674 430
rect 60790 345 61458 430
rect 61574 345 62242 430
rect 62358 345 63026 430
rect 63142 345 63810 430
rect 63926 345 64594 430
rect 64710 345 65378 430
rect 65494 345 66162 430
rect 66278 345 66946 430
rect 67062 345 67730 430
rect 67846 345 68514 430
rect 68630 345 69298 430
rect 69414 345 70082 430
rect 70198 345 70866 430
rect 70982 345 71650 430
rect 71766 345 72434 430
rect 72550 345 73218 430
rect 73334 345 74002 430
rect 74118 345 74786 430
rect 74902 345 75570 430
rect 75686 345 76354 430
rect 76470 345 77138 430
rect 77254 345 77922 430
rect 78038 345 78706 430
rect 78822 345 79490 430
<< metal3 >>
rect 79600 59472 80000 59528
rect 0 59360 400 59416
rect 0 58576 400 58632
rect 79600 58576 80000 58632
rect 0 57792 400 57848
rect 79600 57680 80000 57736
rect 0 57008 400 57064
rect 79600 56784 80000 56840
rect 0 56224 400 56280
rect 79600 55888 80000 55944
rect 0 55440 400 55496
rect 79600 54992 80000 55048
rect 0 54656 400 54712
rect 79600 54096 80000 54152
rect 0 53872 400 53928
rect 79600 53200 80000 53256
rect 0 53088 400 53144
rect 0 52304 400 52360
rect 79600 52304 80000 52360
rect 0 51520 400 51576
rect 79600 51408 80000 51464
rect 0 50736 400 50792
rect 79600 50512 80000 50568
rect 0 49952 400 50008
rect 79600 49616 80000 49672
rect 0 49168 400 49224
rect 79600 48720 80000 48776
rect 0 48384 400 48440
rect 79600 47824 80000 47880
rect 0 47600 400 47656
rect 79600 46928 80000 46984
rect 0 46816 400 46872
rect 0 46032 400 46088
rect 79600 46032 80000 46088
rect 0 45248 400 45304
rect 79600 45136 80000 45192
rect 0 44464 400 44520
rect 79600 44240 80000 44296
rect 0 43680 400 43736
rect 79600 43344 80000 43400
rect 0 42896 400 42952
rect 79600 42448 80000 42504
rect 0 42112 400 42168
rect 79600 41552 80000 41608
rect 0 41328 400 41384
rect 79600 40656 80000 40712
rect 0 40544 400 40600
rect 0 39760 400 39816
rect 79600 39760 80000 39816
rect 0 38976 400 39032
rect 79600 38864 80000 38920
rect 0 38192 400 38248
rect 79600 37968 80000 38024
rect 0 37408 400 37464
rect 79600 37072 80000 37128
rect 0 36624 400 36680
rect 79600 36176 80000 36232
rect 0 35840 400 35896
rect 79600 35280 80000 35336
rect 0 35056 400 35112
rect 79600 34384 80000 34440
rect 0 34272 400 34328
rect 0 33488 400 33544
rect 79600 33488 80000 33544
rect 0 32704 400 32760
rect 79600 32592 80000 32648
rect 0 31920 400 31976
rect 79600 31696 80000 31752
rect 0 31136 400 31192
rect 79600 30800 80000 30856
rect 0 30352 400 30408
rect 79600 29904 80000 29960
rect 0 29568 400 29624
rect 79600 29008 80000 29064
rect 0 28784 400 28840
rect 79600 28112 80000 28168
rect 0 28000 400 28056
rect 0 27216 400 27272
rect 79600 27216 80000 27272
rect 0 26432 400 26488
rect 79600 26320 80000 26376
rect 0 25648 400 25704
rect 79600 25424 80000 25480
rect 0 24864 400 24920
rect 79600 24528 80000 24584
rect 0 24080 400 24136
rect 79600 23632 80000 23688
rect 0 23296 400 23352
rect 79600 22736 80000 22792
rect 0 22512 400 22568
rect 79600 21840 80000 21896
rect 0 21728 400 21784
rect 0 20944 400 21000
rect 79600 20944 80000 21000
rect 0 20160 400 20216
rect 79600 20048 80000 20104
rect 0 19376 400 19432
rect 79600 19152 80000 19208
rect 0 18592 400 18648
rect 79600 18256 80000 18312
rect 0 17808 400 17864
rect 79600 17360 80000 17416
rect 0 17024 400 17080
rect 79600 16464 80000 16520
rect 0 16240 400 16296
rect 79600 15568 80000 15624
rect 0 15456 400 15512
rect 0 14672 400 14728
rect 79600 14672 80000 14728
rect 0 13888 400 13944
rect 79600 13776 80000 13832
rect 0 13104 400 13160
rect 79600 12880 80000 12936
rect 0 12320 400 12376
rect 79600 11984 80000 12040
rect 0 11536 400 11592
rect 79600 11088 80000 11144
rect 0 10752 400 10808
rect 79600 10192 80000 10248
rect 0 9968 400 10024
rect 79600 9296 80000 9352
rect 0 9184 400 9240
rect 0 8400 400 8456
rect 79600 8400 80000 8456
rect 0 7616 400 7672
rect 79600 7504 80000 7560
rect 0 6832 400 6888
rect 79600 6608 80000 6664
rect 0 6048 400 6104
rect 79600 5712 80000 5768
rect 0 5264 400 5320
rect 79600 4816 80000 4872
rect 0 4480 400 4536
rect 79600 3920 80000 3976
rect 0 3696 400 3752
rect 79600 3024 80000 3080
rect 0 2912 400 2968
rect 0 2128 400 2184
rect 79600 2128 80000 2184
rect 0 1344 400 1400
rect 79600 1232 80000 1288
rect 0 560 400 616
rect 79600 336 80000 392
<< obsm3 >>
rect 345 59446 79570 59514
rect 430 59442 79570 59446
rect 430 59330 79674 59442
rect 345 58662 79674 59330
rect 430 58546 79570 58662
rect 345 57878 79674 58546
rect 430 57766 79674 57878
rect 430 57762 79570 57766
rect 345 57650 79570 57762
rect 345 57094 79674 57650
rect 430 56978 79674 57094
rect 345 56870 79674 56978
rect 345 56754 79570 56870
rect 345 56310 79674 56754
rect 430 56194 79674 56310
rect 345 55974 79674 56194
rect 345 55858 79570 55974
rect 345 55526 79674 55858
rect 430 55410 79674 55526
rect 345 55078 79674 55410
rect 345 54962 79570 55078
rect 345 54742 79674 54962
rect 430 54626 79674 54742
rect 345 54182 79674 54626
rect 345 54066 79570 54182
rect 345 53958 79674 54066
rect 430 53842 79674 53958
rect 345 53286 79674 53842
rect 345 53174 79570 53286
rect 430 53170 79570 53174
rect 430 53058 79674 53170
rect 345 52390 79674 53058
rect 430 52274 79570 52390
rect 345 51606 79674 52274
rect 430 51494 79674 51606
rect 430 51490 79570 51494
rect 345 51378 79570 51490
rect 345 50822 79674 51378
rect 430 50706 79674 50822
rect 345 50598 79674 50706
rect 345 50482 79570 50598
rect 345 50038 79674 50482
rect 430 49922 79674 50038
rect 345 49702 79674 49922
rect 345 49586 79570 49702
rect 345 49254 79674 49586
rect 430 49138 79674 49254
rect 345 48806 79674 49138
rect 345 48690 79570 48806
rect 345 48470 79674 48690
rect 430 48354 79674 48470
rect 345 47910 79674 48354
rect 345 47794 79570 47910
rect 345 47686 79674 47794
rect 430 47570 79674 47686
rect 345 47014 79674 47570
rect 345 46902 79570 47014
rect 430 46898 79570 46902
rect 430 46786 79674 46898
rect 345 46118 79674 46786
rect 430 46002 79570 46118
rect 345 45334 79674 46002
rect 430 45222 79674 45334
rect 430 45218 79570 45222
rect 345 45106 79570 45218
rect 345 44550 79674 45106
rect 430 44434 79674 44550
rect 345 44326 79674 44434
rect 345 44210 79570 44326
rect 345 43766 79674 44210
rect 430 43650 79674 43766
rect 345 43430 79674 43650
rect 345 43314 79570 43430
rect 345 42982 79674 43314
rect 430 42866 79674 42982
rect 345 42534 79674 42866
rect 345 42418 79570 42534
rect 345 42198 79674 42418
rect 430 42082 79674 42198
rect 345 41638 79674 42082
rect 345 41522 79570 41638
rect 345 41414 79674 41522
rect 430 41298 79674 41414
rect 345 40742 79674 41298
rect 345 40630 79570 40742
rect 430 40626 79570 40630
rect 430 40514 79674 40626
rect 345 39846 79674 40514
rect 430 39730 79570 39846
rect 345 39062 79674 39730
rect 430 38950 79674 39062
rect 430 38946 79570 38950
rect 345 38834 79570 38946
rect 345 38278 79674 38834
rect 430 38162 79674 38278
rect 345 38054 79674 38162
rect 345 37938 79570 38054
rect 345 37494 79674 37938
rect 430 37378 79674 37494
rect 345 37158 79674 37378
rect 345 37042 79570 37158
rect 345 36710 79674 37042
rect 430 36594 79674 36710
rect 345 36262 79674 36594
rect 345 36146 79570 36262
rect 345 35926 79674 36146
rect 430 35810 79674 35926
rect 345 35366 79674 35810
rect 345 35250 79570 35366
rect 345 35142 79674 35250
rect 430 35026 79674 35142
rect 345 34470 79674 35026
rect 345 34358 79570 34470
rect 430 34354 79570 34358
rect 430 34242 79674 34354
rect 345 33574 79674 34242
rect 430 33458 79570 33574
rect 345 32790 79674 33458
rect 430 32678 79674 32790
rect 430 32674 79570 32678
rect 345 32562 79570 32674
rect 345 32006 79674 32562
rect 430 31890 79674 32006
rect 345 31782 79674 31890
rect 345 31666 79570 31782
rect 345 31222 79674 31666
rect 430 31106 79674 31222
rect 345 30886 79674 31106
rect 345 30770 79570 30886
rect 345 30438 79674 30770
rect 430 30322 79674 30438
rect 345 29990 79674 30322
rect 345 29874 79570 29990
rect 345 29654 79674 29874
rect 430 29538 79674 29654
rect 345 29094 79674 29538
rect 345 28978 79570 29094
rect 345 28870 79674 28978
rect 430 28754 79674 28870
rect 345 28198 79674 28754
rect 345 28086 79570 28198
rect 430 28082 79570 28086
rect 430 27970 79674 28082
rect 345 27302 79674 27970
rect 430 27186 79570 27302
rect 345 26518 79674 27186
rect 430 26406 79674 26518
rect 430 26402 79570 26406
rect 345 26290 79570 26402
rect 345 25734 79674 26290
rect 430 25618 79674 25734
rect 345 25510 79674 25618
rect 345 25394 79570 25510
rect 345 24950 79674 25394
rect 430 24834 79674 24950
rect 345 24614 79674 24834
rect 345 24498 79570 24614
rect 345 24166 79674 24498
rect 430 24050 79674 24166
rect 345 23718 79674 24050
rect 345 23602 79570 23718
rect 345 23382 79674 23602
rect 430 23266 79674 23382
rect 345 22822 79674 23266
rect 345 22706 79570 22822
rect 345 22598 79674 22706
rect 430 22482 79674 22598
rect 345 21926 79674 22482
rect 345 21814 79570 21926
rect 430 21810 79570 21814
rect 430 21698 79674 21810
rect 345 21030 79674 21698
rect 430 20914 79570 21030
rect 345 20246 79674 20914
rect 430 20134 79674 20246
rect 430 20130 79570 20134
rect 345 20018 79570 20130
rect 345 19462 79674 20018
rect 430 19346 79674 19462
rect 345 19238 79674 19346
rect 345 19122 79570 19238
rect 345 18678 79674 19122
rect 430 18562 79674 18678
rect 345 18342 79674 18562
rect 345 18226 79570 18342
rect 345 17894 79674 18226
rect 430 17778 79674 17894
rect 345 17446 79674 17778
rect 345 17330 79570 17446
rect 345 17110 79674 17330
rect 430 16994 79674 17110
rect 345 16550 79674 16994
rect 345 16434 79570 16550
rect 345 16326 79674 16434
rect 430 16210 79674 16326
rect 345 15654 79674 16210
rect 345 15542 79570 15654
rect 430 15538 79570 15542
rect 430 15426 79674 15538
rect 345 14758 79674 15426
rect 430 14642 79570 14758
rect 345 13974 79674 14642
rect 430 13862 79674 13974
rect 430 13858 79570 13862
rect 345 13746 79570 13858
rect 345 13190 79674 13746
rect 430 13074 79674 13190
rect 345 12966 79674 13074
rect 345 12850 79570 12966
rect 345 12406 79674 12850
rect 430 12290 79674 12406
rect 345 12070 79674 12290
rect 345 11954 79570 12070
rect 345 11622 79674 11954
rect 430 11506 79674 11622
rect 345 11174 79674 11506
rect 345 11058 79570 11174
rect 345 10838 79674 11058
rect 430 10722 79674 10838
rect 345 10278 79674 10722
rect 345 10162 79570 10278
rect 345 10054 79674 10162
rect 430 9938 79674 10054
rect 345 9382 79674 9938
rect 345 9270 79570 9382
rect 430 9266 79570 9270
rect 430 9154 79674 9266
rect 345 8486 79674 9154
rect 430 8370 79570 8486
rect 345 7702 79674 8370
rect 430 7590 79674 7702
rect 430 7586 79570 7590
rect 345 7474 79570 7586
rect 345 6918 79674 7474
rect 430 6802 79674 6918
rect 345 6694 79674 6802
rect 345 6578 79570 6694
rect 345 6134 79674 6578
rect 430 6018 79674 6134
rect 345 5798 79674 6018
rect 345 5682 79570 5798
rect 345 5350 79674 5682
rect 430 5234 79674 5350
rect 345 4902 79674 5234
rect 345 4786 79570 4902
rect 345 4566 79674 4786
rect 430 4450 79674 4566
rect 345 4006 79674 4450
rect 345 3890 79570 4006
rect 345 3782 79674 3890
rect 430 3666 79674 3782
rect 345 3110 79674 3666
rect 345 2998 79570 3110
rect 430 2994 79570 2998
rect 430 2882 79674 2994
rect 345 2214 79674 2882
rect 430 2098 79570 2214
rect 345 1430 79674 2098
rect 430 1318 79674 1430
rect 430 1314 79570 1318
rect 345 1202 79570 1314
rect 345 646 79674 1202
rect 430 530 79674 646
rect 345 422 79674 530
rect 345 350 79570 422
<< metal4 >>
rect 2224 1538 2384 58438
rect 9904 1538 10064 58438
rect 17584 1538 17744 58438
rect 25264 1538 25424 58438
rect 32944 1538 33104 58438
rect 40624 1538 40784 58438
rect 48304 1538 48464 58438
rect 55984 1538 56144 58438
rect 63664 1538 63824 58438
rect 71344 1538 71504 58438
rect 79024 1538 79184 58438
<< obsm4 >>
rect 5502 2137 9874 58343
rect 10094 2137 17554 58343
rect 17774 2137 25234 58343
rect 25454 2137 32914 58343
rect 33134 2137 40594 58343
rect 40814 2137 48274 58343
rect 48494 2137 55954 58343
rect 56174 2137 63634 58343
rect 63854 2137 71314 58343
rect 71534 2137 78610 58343
<< labels >>
rlabel metal2 s 2576 59600 2632 60000 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 22736 59600 22792 60000 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 24752 59600 24808 60000 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 26768 59600 26824 60000 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 28784 59600 28840 60000 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 30800 59600 30856 60000 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 32816 59600 32872 60000 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 34832 59600 34888 60000 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 36848 59600 36904 60000 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 38864 59600 38920 60000 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 40880 59600 40936 60000 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 4592 59600 4648 60000 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 42896 59600 42952 60000 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 44912 59600 44968 60000 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 46928 59600 46984 60000 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 48944 59600 49000 60000 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 50960 59600 51016 60000 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 52976 59600 53032 60000 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 54992 59600 55048 60000 6 io_in[26]
port 19 nsew signal input
rlabel metal2 s 57008 59600 57064 60000 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 59024 59600 59080 60000 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 61040 59600 61096 60000 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 6608 59600 6664 60000 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 63056 59600 63112 60000 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 65072 59600 65128 60000 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 67088 59600 67144 60000 6 io_in[32]
port 26 nsew signal input
rlabel metal2 s 69104 59600 69160 60000 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 71120 59600 71176 60000 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 73136 59600 73192 60000 6 io_in[35]
port 29 nsew signal input
rlabel metal2 s 75152 59600 75208 60000 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 77168 59600 77224 60000 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 8624 59600 8680 60000 6 io_in[3]
port 32 nsew signal input
rlabel metal2 s 10640 59600 10696 60000 6 io_in[4]
port 33 nsew signal input
rlabel metal2 s 12656 59600 12712 60000 6 io_in[5]
port 34 nsew signal input
rlabel metal2 s 14672 59600 14728 60000 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 16688 59600 16744 60000 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 18704 59600 18760 60000 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 20720 59600 20776 60000 6 io_in[9]
port 38 nsew signal input
rlabel metal3 s 0 30352 400 30408 6 io_oeb[0]
port 39 nsew signal output
rlabel metal3 s 0 38192 400 38248 6 io_oeb[10]
port 40 nsew signal output
rlabel metal3 s 0 38976 400 39032 6 io_oeb[11]
port 41 nsew signal output
rlabel metal3 s 0 39760 400 39816 6 io_oeb[12]
port 42 nsew signal output
rlabel metal3 s 0 40544 400 40600 6 io_oeb[13]
port 43 nsew signal output
rlabel metal3 s 0 41328 400 41384 6 io_oeb[14]
port 44 nsew signal output
rlabel metal3 s 0 42112 400 42168 6 io_oeb[15]
port 45 nsew signal output
rlabel metal3 s 0 42896 400 42952 6 io_oeb[16]
port 46 nsew signal output
rlabel metal3 s 0 43680 400 43736 6 io_oeb[17]
port 47 nsew signal output
rlabel metal3 s 0 44464 400 44520 6 io_oeb[18]
port 48 nsew signal output
rlabel metal3 s 0 45248 400 45304 6 io_oeb[19]
port 49 nsew signal output
rlabel metal3 s 0 31136 400 31192 6 io_oeb[1]
port 50 nsew signal output
rlabel metal3 s 0 46032 400 46088 6 io_oeb[20]
port 51 nsew signal output
rlabel metal3 s 0 46816 400 46872 6 io_oeb[21]
port 52 nsew signal output
rlabel metal3 s 0 47600 400 47656 6 io_oeb[22]
port 53 nsew signal output
rlabel metal3 s 0 48384 400 48440 6 io_oeb[23]
port 54 nsew signal output
rlabel metal3 s 0 49168 400 49224 6 io_oeb[24]
port 55 nsew signal output
rlabel metal3 s 0 49952 400 50008 6 io_oeb[25]
port 56 nsew signal output
rlabel metal3 s 0 50736 400 50792 6 io_oeb[26]
port 57 nsew signal output
rlabel metal3 s 0 51520 400 51576 6 io_oeb[27]
port 58 nsew signal output
rlabel metal3 s 0 52304 400 52360 6 io_oeb[28]
port 59 nsew signal output
rlabel metal3 s 0 53088 400 53144 6 io_oeb[29]
port 60 nsew signal output
rlabel metal3 s 0 31920 400 31976 6 io_oeb[2]
port 61 nsew signal output
rlabel metal3 s 0 53872 400 53928 6 io_oeb[30]
port 62 nsew signal output
rlabel metal3 s 0 54656 400 54712 6 io_oeb[31]
port 63 nsew signal output
rlabel metal3 s 0 55440 400 55496 6 io_oeb[32]
port 64 nsew signal output
rlabel metal3 s 0 56224 400 56280 6 io_oeb[33]
port 65 nsew signal output
rlabel metal3 s 0 57008 400 57064 6 io_oeb[34]
port 66 nsew signal output
rlabel metal3 s 0 57792 400 57848 6 io_oeb[35]
port 67 nsew signal output
rlabel metal3 s 0 58576 400 58632 6 io_oeb[36]
port 68 nsew signal output
rlabel metal3 s 0 59360 400 59416 6 io_oeb[37]
port 69 nsew signal output
rlabel metal3 s 0 32704 400 32760 6 io_oeb[3]
port 70 nsew signal output
rlabel metal3 s 0 33488 400 33544 6 io_oeb[4]
port 71 nsew signal output
rlabel metal3 s 0 34272 400 34328 6 io_oeb[5]
port 72 nsew signal output
rlabel metal3 s 0 35056 400 35112 6 io_oeb[6]
port 73 nsew signal output
rlabel metal3 s 0 35840 400 35896 6 io_oeb[7]
port 74 nsew signal output
rlabel metal3 s 0 36624 400 36680 6 io_oeb[8]
port 75 nsew signal output
rlabel metal3 s 0 37408 400 37464 6 io_oeb[9]
port 76 nsew signal output
rlabel metal3 s 0 560 400 616 6 io_out[0]
port 77 nsew signal output
rlabel metal3 s 0 8400 400 8456 6 io_out[10]
port 78 nsew signal output
rlabel metal3 s 0 9184 400 9240 6 io_out[11]
port 79 nsew signal output
rlabel metal3 s 0 9968 400 10024 6 io_out[12]
port 80 nsew signal output
rlabel metal3 s 0 10752 400 10808 6 io_out[13]
port 81 nsew signal output
rlabel metal3 s 0 11536 400 11592 6 io_out[14]
port 82 nsew signal output
rlabel metal3 s 0 12320 400 12376 6 io_out[15]
port 83 nsew signal output
rlabel metal3 s 0 13104 400 13160 6 io_out[16]
port 84 nsew signal output
rlabel metal3 s 0 13888 400 13944 6 io_out[17]
port 85 nsew signal output
rlabel metal3 s 0 14672 400 14728 6 io_out[18]
port 86 nsew signal output
rlabel metal3 s 0 15456 400 15512 6 io_out[19]
port 87 nsew signal output
rlabel metal3 s 0 1344 400 1400 6 io_out[1]
port 88 nsew signal output
rlabel metal3 s 0 16240 400 16296 6 io_out[20]
port 89 nsew signal output
rlabel metal3 s 0 17024 400 17080 6 io_out[21]
port 90 nsew signal output
rlabel metal3 s 0 17808 400 17864 6 io_out[22]
port 91 nsew signal output
rlabel metal3 s 0 18592 400 18648 6 io_out[23]
port 92 nsew signal output
rlabel metal3 s 0 19376 400 19432 6 io_out[24]
port 93 nsew signal output
rlabel metal3 s 0 20160 400 20216 6 io_out[25]
port 94 nsew signal output
rlabel metal3 s 0 20944 400 21000 6 io_out[26]
port 95 nsew signal output
rlabel metal3 s 0 21728 400 21784 6 io_out[27]
port 96 nsew signal output
rlabel metal3 s 0 22512 400 22568 6 io_out[28]
port 97 nsew signal output
rlabel metal3 s 0 23296 400 23352 6 io_out[29]
port 98 nsew signal output
rlabel metal3 s 0 2128 400 2184 6 io_out[2]
port 99 nsew signal output
rlabel metal3 s 0 24080 400 24136 6 io_out[30]
port 100 nsew signal output
rlabel metal3 s 0 24864 400 24920 6 io_out[31]
port 101 nsew signal output
rlabel metal3 s 0 25648 400 25704 6 io_out[32]
port 102 nsew signal output
rlabel metal3 s 0 26432 400 26488 6 io_out[33]
port 103 nsew signal output
rlabel metal3 s 0 27216 400 27272 6 io_out[34]
port 104 nsew signal output
rlabel metal3 s 0 28000 400 28056 6 io_out[35]
port 105 nsew signal output
rlabel metal3 s 0 28784 400 28840 6 io_out[36]
port 106 nsew signal output
rlabel metal3 s 0 29568 400 29624 6 io_out[37]
port 107 nsew signal output
rlabel metal3 s 0 2912 400 2968 6 io_out[3]
port 108 nsew signal output
rlabel metal3 s 0 3696 400 3752 6 io_out[4]
port 109 nsew signal output
rlabel metal3 s 0 4480 400 4536 6 io_out[5]
port 110 nsew signal output
rlabel metal3 s 0 5264 400 5320 6 io_out[6]
port 111 nsew signal output
rlabel metal3 s 0 6048 400 6104 6 io_out[7]
port 112 nsew signal output
rlabel metal3 s 0 6832 400 6888 6 io_out[8]
port 113 nsew signal output
rlabel metal3 s 0 7616 400 7672 6 io_out[9]
port 114 nsew signal output
rlabel metal3 s 79600 57680 80000 57736 6 irq[0]
port 115 nsew signal output
rlabel metal3 s 79600 58576 80000 58632 6 irq[1]
port 116 nsew signal output
rlabel metal3 s 79600 59472 80000 59528 6 irq[2]
port 117 nsew signal output
rlabel metal3 s 79600 336 80000 392 6 la_data_out[0]
port 118 nsew signal output
rlabel metal3 s 79600 9296 80000 9352 6 la_data_out[10]
port 119 nsew signal output
rlabel metal3 s 79600 10192 80000 10248 6 la_data_out[11]
port 120 nsew signal output
rlabel metal3 s 79600 11088 80000 11144 6 la_data_out[12]
port 121 nsew signal output
rlabel metal3 s 79600 11984 80000 12040 6 la_data_out[13]
port 122 nsew signal output
rlabel metal3 s 79600 12880 80000 12936 6 la_data_out[14]
port 123 nsew signal output
rlabel metal3 s 79600 13776 80000 13832 6 la_data_out[15]
port 124 nsew signal output
rlabel metal3 s 79600 14672 80000 14728 6 la_data_out[16]
port 125 nsew signal output
rlabel metal3 s 79600 15568 80000 15624 6 la_data_out[17]
port 126 nsew signal output
rlabel metal3 s 79600 16464 80000 16520 6 la_data_out[18]
port 127 nsew signal output
rlabel metal3 s 79600 17360 80000 17416 6 la_data_out[19]
port 128 nsew signal output
rlabel metal3 s 79600 1232 80000 1288 6 la_data_out[1]
port 129 nsew signal output
rlabel metal3 s 79600 18256 80000 18312 6 la_data_out[20]
port 130 nsew signal output
rlabel metal3 s 79600 19152 80000 19208 6 la_data_out[21]
port 131 nsew signal output
rlabel metal3 s 79600 20048 80000 20104 6 la_data_out[22]
port 132 nsew signal output
rlabel metal3 s 79600 20944 80000 21000 6 la_data_out[23]
port 133 nsew signal output
rlabel metal3 s 79600 21840 80000 21896 6 la_data_out[24]
port 134 nsew signal output
rlabel metal3 s 79600 22736 80000 22792 6 la_data_out[25]
port 135 nsew signal output
rlabel metal3 s 79600 23632 80000 23688 6 la_data_out[26]
port 136 nsew signal output
rlabel metal3 s 79600 24528 80000 24584 6 la_data_out[27]
port 137 nsew signal output
rlabel metal3 s 79600 25424 80000 25480 6 la_data_out[28]
port 138 nsew signal output
rlabel metal3 s 79600 26320 80000 26376 6 la_data_out[29]
port 139 nsew signal output
rlabel metal3 s 79600 2128 80000 2184 6 la_data_out[2]
port 140 nsew signal output
rlabel metal3 s 79600 27216 80000 27272 6 la_data_out[30]
port 141 nsew signal output
rlabel metal3 s 79600 28112 80000 28168 6 la_data_out[31]
port 142 nsew signal output
rlabel metal3 s 79600 29008 80000 29064 6 la_data_out[32]
port 143 nsew signal output
rlabel metal3 s 79600 29904 80000 29960 6 la_data_out[33]
port 144 nsew signal output
rlabel metal3 s 79600 30800 80000 30856 6 la_data_out[34]
port 145 nsew signal output
rlabel metal3 s 79600 31696 80000 31752 6 la_data_out[35]
port 146 nsew signal output
rlabel metal3 s 79600 32592 80000 32648 6 la_data_out[36]
port 147 nsew signal output
rlabel metal3 s 79600 33488 80000 33544 6 la_data_out[37]
port 148 nsew signal output
rlabel metal3 s 79600 34384 80000 34440 6 la_data_out[38]
port 149 nsew signal output
rlabel metal3 s 79600 35280 80000 35336 6 la_data_out[39]
port 150 nsew signal output
rlabel metal3 s 79600 3024 80000 3080 6 la_data_out[3]
port 151 nsew signal output
rlabel metal3 s 79600 36176 80000 36232 6 la_data_out[40]
port 152 nsew signal output
rlabel metal3 s 79600 37072 80000 37128 6 la_data_out[41]
port 153 nsew signal output
rlabel metal3 s 79600 37968 80000 38024 6 la_data_out[42]
port 154 nsew signal output
rlabel metal3 s 79600 38864 80000 38920 6 la_data_out[43]
port 155 nsew signal output
rlabel metal3 s 79600 39760 80000 39816 6 la_data_out[44]
port 156 nsew signal output
rlabel metal3 s 79600 40656 80000 40712 6 la_data_out[45]
port 157 nsew signal output
rlabel metal3 s 79600 41552 80000 41608 6 la_data_out[46]
port 158 nsew signal output
rlabel metal3 s 79600 42448 80000 42504 6 la_data_out[47]
port 159 nsew signal output
rlabel metal3 s 79600 43344 80000 43400 6 la_data_out[48]
port 160 nsew signal output
rlabel metal3 s 79600 44240 80000 44296 6 la_data_out[49]
port 161 nsew signal output
rlabel metal3 s 79600 3920 80000 3976 6 la_data_out[4]
port 162 nsew signal output
rlabel metal3 s 79600 45136 80000 45192 6 la_data_out[50]
port 163 nsew signal output
rlabel metal3 s 79600 46032 80000 46088 6 la_data_out[51]
port 164 nsew signal output
rlabel metal3 s 79600 46928 80000 46984 6 la_data_out[52]
port 165 nsew signal output
rlabel metal3 s 79600 47824 80000 47880 6 la_data_out[53]
port 166 nsew signal output
rlabel metal3 s 79600 48720 80000 48776 6 la_data_out[54]
port 167 nsew signal output
rlabel metal3 s 79600 49616 80000 49672 6 la_data_out[55]
port 168 nsew signal output
rlabel metal3 s 79600 50512 80000 50568 6 la_data_out[56]
port 169 nsew signal output
rlabel metal3 s 79600 51408 80000 51464 6 la_data_out[57]
port 170 nsew signal output
rlabel metal3 s 79600 52304 80000 52360 6 la_data_out[58]
port 171 nsew signal output
rlabel metal3 s 79600 53200 80000 53256 6 la_data_out[59]
port 172 nsew signal output
rlabel metal3 s 79600 4816 80000 4872 6 la_data_out[5]
port 173 nsew signal output
rlabel metal3 s 79600 54096 80000 54152 6 la_data_out[60]
port 174 nsew signal output
rlabel metal3 s 79600 54992 80000 55048 6 la_data_out[61]
port 175 nsew signal output
rlabel metal3 s 79600 55888 80000 55944 6 la_data_out[62]
port 176 nsew signal output
rlabel metal3 s 79600 56784 80000 56840 6 la_data_out[63]
port 177 nsew signal output
rlabel metal3 s 79600 5712 80000 5768 6 la_data_out[6]
port 178 nsew signal output
rlabel metal3 s 79600 6608 80000 6664 6 la_data_out[7]
port 179 nsew signal output
rlabel metal3 s 79600 7504 80000 7560 6 la_data_out[8]
port 180 nsew signal output
rlabel metal3 s 79600 8400 80000 8456 6 la_data_out[9]
port 181 nsew signal output
rlabel metal4 s 2224 1538 2384 58438 6 vdd
port 182 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 58438 6 vdd
port 182 nsew power bidirectional
rlabel metal4 s 32944 1538 33104 58438 6 vdd
port 182 nsew power bidirectional
rlabel metal4 s 48304 1538 48464 58438 6 vdd
port 182 nsew power bidirectional
rlabel metal4 s 63664 1538 63824 58438 6 vdd
port 182 nsew power bidirectional
rlabel metal4 s 79024 1538 79184 58438 6 vdd
port 182 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 58438 6 vss
port 183 nsew ground bidirectional
rlabel metal4 s 25264 1538 25424 58438 6 vss
port 183 nsew ground bidirectional
rlabel metal4 s 40624 1538 40784 58438 6 vss
port 183 nsew ground bidirectional
rlabel metal4 s 55984 1538 56144 58438 6 vss
port 183 nsew ground bidirectional
rlabel metal4 s 71344 1538 71504 58438 6 vss
port 183 nsew ground bidirectional
rlabel metal2 s 336 0 392 400 6 wb_clk_i
port 184 nsew signal input
rlabel metal2 s 1120 0 1176 400 6 wb_rst_i
port 185 nsew signal input
rlabel metal2 s 1904 0 1960 400 6 wbs_ack_o
port 186 nsew signal output
rlabel metal2 s 5040 0 5096 400 6 wbs_adr_i[0]
port 187 nsew signal input
rlabel metal2 s 28560 0 28616 400 6 wbs_adr_i[10]
port 188 nsew signal input
rlabel metal2 s 30912 0 30968 400 6 wbs_adr_i[11]
port 189 nsew signal input
rlabel metal2 s 33264 0 33320 400 6 wbs_adr_i[12]
port 190 nsew signal input
rlabel metal2 s 35616 0 35672 400 6 wbs_adr_i[13]
port 191 nsew signal input
rlabel metal2 s 37968 0 38024 400 6 wbs_adr_i[14]
port 192 nsew signal input
rlabel metal2 s 40320 0 40376 400 6 wbs_adr_i[15]
port 193 nsew signal input
rlabel metal2 s 42672 0 42728 400 6 wbs_adr_i[16]
port 194 nsew signal input
rlabel metal2 s 45024 0 45080 400 6 wbs_adr_i[17]
port 195 nsew signal input
rlabel metal2 s 47376 0 47432 400 6 wbs_adr_i[18]
port 196 nsew signal input
rlabel metal2 s 49728 0 49784 400 6 wbs_adr_i[19]
port 197 nsew signal input
rlabel metal2 s 7392 0 7448 400 6 wbs_adr_i[1]
port 198 nsew signal input
rlabel metal2 s 52080 0 52136 400 6 wbs_adr_i[20]
port 199 nsew signal input
rlabel metal2 s 54432 0 54488 400 6 wbs_adr_i[21]
port 200 nsew signal input
rlabel metal2 s 56784 0 56840 400 6 wbs_adr_i[22]
port 201 nsew signal input
rlabel metal2 s 59136 0 59192 400 6 wbs_adr_i[23]
port 202 nsew signal input
rlabel metal2 s 61488 0 61544 400 6 wbs_adr_i[24]
port 203 nsew signal input
rlabel metal2 s 63840 0 63896 400 6 wbs_adr_i[25]
port 204 nsew signal input
rlabel metal2 s 66192 0 66248 400 6 wbs_adr_i[26]
port 205 nsew signal input
rlabel metal2 s 68544 0 68600 400 6 wbs_adr_i[27]
port 206 nsew signal input
rlabel metal2 s 70896 0 70952 400 6 wbs_adr_i[28]
port 207 nsew signal input
rlabel metal2 s 73248 0 73304 400 6 wbs_adr_i[29]
port 208 nsew signal input
rlabel metal2 s 9744 0 9800 400 6 wbs_adr_i[2]
port 209 nsew signal input
rlabel metal2 s 75600 0 75656 400 6 wbs_adr_i[30]
port 210 nsew signal input
rlabel metal2 s 77952 0 78008 400 6 wbs_adr_i[31]
port 211 nsew signal input
rlabel metal2 s 12096 0 12152 400 6 wbs_adr_i[3]
port 212 nsew signal input
rlabel metal2 s 14448 0 14504 400 6 wbs_adr_i[4]
port 213 nsew signal input
rlabel metal2 s 16800 0 16856 400 6 wbs_adr_i[5]
port 214 nsew signal input
rlabel metal2 s 19152 0 19208 400 6 wbs_adr_i[6]
port 215 nsew signal input
rlabel metal2 s 21504 0 21560 400 6 wbs_adr_i[7]
port 216 nsew signal input
rlabel metal2 s 23856 0 23912 400 6 wbs_adr_i[8]
port 217 nsew signal input
rlabel metal2 s 26208 0 26264 400 6 wbs_adr_i[9]
port 218 nsew signal input
rlabel metal2 s 2688 0 2744 400 6 wbs_cyc_i
port 219 nsew signal input
rlabel metal2 s 5824 0 5880 400 6 wbs_dat_i[0]
port 220 nsew signal input
rlabel metal2 s 29344 0 29400 400 6 wbs_dat_i[10]
port 221 nsew signal input
rlabel metal2 s 31696 0 31752 400 6 wbs_dat_i[11]
port 222 nsew signal input
rlabel metal2 s 34048 0 34104 400 6 wbs_dat_i[12]
port 223 nsew signal input
rlabel metal2 s 36400 0 36456 400 6 wbs_dat_i[13]
port 224 nsew signal input
rlabel metal2 s 38752 0 38808 400 6 wbs_dat_i[14]
port 225 nsew signal input
rlabel metal2 s 41104 0 41160 400 6 wbs_dat_i[15]
port 226 nsew signal input
rlabel metal2 s 43456 0 43512 400 6 wbs_dat_i[16]
port 227 nsew signal input
rlabel metal2 s 45808 0 45864 400 6 wbs_dat_i[17]
port 228 nsew signal input
rlabel metal2 s 48160 0 48216 400 6 wbs_dat_i[18]
port 229 nsew signal input
rlabel metal2 s 50512 0 50568 400 6 wbs_dat_i[19]
port 230 nsew signal input
rlabel metal2 s 8176 0 8232 400 6 wbs_dat_i[1]
port 231 nsew signal input
rlabel metal2 s 52864 0 52920 400 6 wbs_dat_i[20]
port 232 nsew signal input
rlabel metal2 s 55216 0 55272 400 6 wbs_dat_i[21]
port 233 nsew signal input
rlabel metal2 s 57568 0 57624 400 6 wbs_dat_i[22]
port 234 nsew signal input
rlabel metal2 s 59920 0 59976 400 6 wbs_dat_i[23]
port 235 nsew signal input
rlabel metal2 s 62272 0 62328 400 6 wbs_dat_i[24]
port 236 nsew signal input
rlabel metal2 s 64624 0 64680 400 6 wbs_dat_i[25]
port 237 nsew signal input
rlabel metal2 s 66976 0 67032 400 6 wbs_dat_i[26]
port 238 nsew signal input
rlabel metal2 s 69328 0 69384 400 6 wbs_dat_i[27]
port 239 nsew signal input
rlabel metal2 s 71680 0 71736 400 6 wbs_dat_i[28]
port 240 nsew signal input
rlabel metal2 s 74032 0 74088 400 6 wbs_dat_i[29]
port 241 nsew signal input
rlabel metal2 s 10528 0 10584 400 6 wbs_dat_i[2]
port 242 nsew signal input
rlabel metal2 s 76384 0 76440 400 6 wbs_dat_i[30]
port 243 nsew signal input
rlabel metal2 s 78736 0 78792 400 6 wbs_dat_i[31]
port 244 nsew signal input
rlabel metal2 s 12880 0 12936 400 6 wbs_dat_i[3]
port 245 nsew signal input
rlabel metal2 s 15232 0 15288 400 6 wbs_dat_i[4]
port 246 nsew signal input
rlabel metal2 s 17584 0 17640 400 6 wbs_dat_i[5]
port 247 nsew signal input
rlabel metal2 s 19936 0 19992 400 6 wbs_dat_i[6]
port 248 nsew signal input
rlabel metal2 s 22288 0 22344 400 6 wbs_dat_i[7]
port 249 nsew signal input
rlabel metal2 s 24640 0 24696 400 6 wbs_dat_i[8]
port 250 nsew signal input
rlabel metal2 s 26992 0 27048 400 6 wbs_dat_i[9]
port 251 nsew signal input
rlabel metal2 s 6608 0 6664 400 6 wbs_dat_o[0]
port 252 nsew signal output
rlabel metal2 s 30128 0 30184 400 6 wbs_dat_o[10]
port 253 nsew signal output
rlabel metal2 s 32480 0 32536 400 6 wbs_dat_o[11]
port 254 nsew signal output
rlabel metal2 s 34832 0 34888 400 6 wbs_dat_o[12]
port 255 nsew signal output
rlabel metal2 s 37184 0 37240 400 6 wbs_dat_o[13]
port 256 nsew signal output
rlabel metal2 s 39536 0 39592 400 6 wbs_dat_o[14]
port 257 nsew signal output
rlabel metal2 s 41888 0 41944 400 6 wbs_dat_o[15]
port 258 nsew signal output
rlabel metal2 s 44240 0 44296 400 6 wbs_dat_o[16]
port 259 nsew signal output
rlabel metal2 s 46592 0 46648 400 6 wbs_dat_o[17]
port 260 nsew signal output
rlabel metal2 s 48944 0 49000 400 6 wbs_dat_o[18]
port 261 nsew signal output
rlabel metal2 s 51296 0 51352 400 6 wbs_dat_o[19]
port 262 nsew signal output
rlabel metal2 s 8960 0 9016 400 6 wbs_dat_o[1]
port 263 nsew signal output
rlabel metal2 s 53648 0 53704 400 6 wbs_dat_o[20]
port 264 nsew signal output
rlabel metal2 s 56000 0 56056 400 6 wbs_dat_o[21]
port 265 nsew signal output
rlabel metal2 s 58352 0 58408 400 6 wbs_dat_o[22]
port 266 nsew signal output
rlabel metal2 s 60704 0 60760 400 6 wbs_dat_o[23]
port 267 nsew signal output
rlabel metal2 s 63056 0 63112 400 6 wbs_dat_o[24]
port 268 nsew signal output
rlabel metal2 s 65408 0 65464 400 6 wbs_dat_o[25]
port 269 nsew signal output
rlabel metal2 s 67760 0 67816 400 6 wbs_dat_o[26]
port 270 nsew signal output
rlabel metal2 s 70112 0 70168 400 6 wbs_dat_o[27]
port 271 nsew signal output
rlabel metal2 s 72464 0 72520 400 6 wbs_dat_o[28]
port 272 nsew signal output
rlabel metal2 s 74816 0 74872 400 6 wbs_dat_o[29]
port 273 nsew signal output
rlabel metal2 s 11312 0 11368 400 6 wbs_dat_o[2]
port 274 nsew signal output
rlabel metal2 s 77168 0 77224 400 6 wbs_dat_o[30]
port 275 nsew signal output
rlabel metal2 s 79520 0 79576 400 6 wbs_dat_o[31]
port 276 nsew signal output
rlabel metal2 s 13664 0 13720 400 6 wbs_dat_o[3]
port 277 nsew signal output
rlabel metal2 s 16016 0 16072 400 6 wbs_dat_o[4]
port 278 nsew signal output
rlabel metal2 s 18368 0 18424 400 6 wbs_dat_o[5]
port 279 nsew signal output
rlabel metal2 s 20720 0 20776 400 6 wbs_dat_o[6]
port 280 nsew signal output
rlabel metal2 s 23072 0 23128 400 6 wbs_dat_o[7]
port 281 nsew signal output
rlabel metal2 s 25424 0 25480 400 6 wbs_dat_o[8]
port 282 nsew signal output
rlabel metal2 s 27776 0 27832 400 6 wbs_dat_o[9]
port 283 nsew signal output
rlabel metal2 s 3472 0 3528 400 6 wbs_stb_i
port 284 nsew signal input
rlabel metal2 s 4256 0 4312 400 6 wbs_we_i
port 285 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 80000 60000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 12711336
string GDS_FILE /media/lucah/fbc90f8f-67e9-406d-9872-54f02ad6a2d8/AS2650/openlane/wrapped_as2650/runs/23_11_15_15_16/results/signoff/wrapped_as2650.magic.gds
string GDS_START 576422
<< end >>

