magic
tech gf180mcuD
magscale 1 5
timestamp 1700512880
<< obsm1 >>
rect 672 1538 24304 23225
<< metal2 >>
rect 1344 24600 1400 25000
rect 2016 24600 2072 25000
rect 2688 24600 2744 25000
rect 3360 24600 3416 25000
rect 4032 24600 4088 25000
rect 4704 24600 4760 25000
rect 5376 24600 5432 25000
rect 6048 24600 6104 25000
rect 6720 24600 6776 25000
rect 7392 24600 7448 25000
rect 8064 24600 8120 25000
rect 8736 24600 8792 25000
rect 9408 24600 9464 25000
rect 10080 24600 10136 25000
rect 10752 24600 10808 25000
rect 11424 24600 11480 25000
rect 12096 24600 12152 25000
rect 12768 24600 12824 25000
rect 13440 24600 13496 25000
rect 14112 24600 14168 25000
rect 14784 24600 14840 25000
rect 15456 24600 15512 25000
rect 16128 24600 16184 25000
rect 16800 24600 16856 25000
rect 17472 24600 17528 25000
rect 18144 24600 18200 25000
rect 18816 24600 18872 25000
rect 19488 24600 19544 25000
rect 20160 24600 20216 25000
rect 20832 24600 20888 25000
rect 21504 24600 21560 25000
rect 22176 24600 22232 25000
rect 22848 24600 22904 25000
rect 23520 24600 23576 25000
rect 1344 0 1400 400
rect 2352 0 2408 400
rect 3360 0 3416 400
rect 4368 0 4424 400
rect 5376 0 5432 400
rect 6384 0 6440 400
rect 7392 0 7448 400
rect 8400 0 8456 400
rect 9408 0 9464 400
rect 10416 0 10472 400
rect 11424 0 11480 400
rect 12432 0 12488 400
rect 13440 0 13496 400
rect 14448 0 14504 400
rect 15456 0 15512 400
rect 16464 0 16520 400
rect 17472 0 17528 400
rect 18480 0 18536 400
rect 19488 0 19544 400
rect 20496 0 20552 400
rect 21504 0 21560 400
rect 22512 0 22568 400
rect 23520 0 23576 400
<< obsm2 >>
rect 742 24570 1314 24682
rect 1430 24570 1986 24682
rect 2102 24570 2658 24682
rect 2774 24570 3330 24682
rect 3446 24570 4002 24682
rect 4118 24570 4674 24682
rect 4790 24570 5346 24682
rect 5462 24570 6018 24682
rect 6134 24570 6690 24682
rect 6806 24570 7362 24682
rect 7478 24570 8034 24682
rect 8150 24570 8706 24682
rect 8822 24570 9378 24682
rect 9494 24570 10050 24682
rect 10166 24570 10722 24682
rect 10838 24570 11394 24682
rect 11510 24570 12066 24682
rect 12182 24570 12738 24682
rect 12854 24570 13410 24682
rect 13526 24570 14082 24682
rect 14198 24570 14754 24682
rect 14870 24570 15426 24682
rect 15542 24570 16098 24682
rect 16214 24570 16770 24682
rect 16886 24570 17442 24682
rect 17558 24570 18114 24682
rect 18230 24570 18786 24682
rect 18902 24570 19458 24682
rect 19574 24570 20130 24682
rect 20246 24570 20802 24682
rect 20918 24570 21474 24682
rect 21590 24570 22146 24682
rect 22262 24570 22818 24682
rect 22934 24570 23490 24682
rect 23606 24570 24122 24682
rect 742 430 24122 24570
rect 742 400 1314 430
rect 1430 400 2322 430
rect 2438 400 3330 430
rect 3446 400 4338 430
rect 4454 400 5346 430
rect 5462 400 6354 430
rect 6470 400 7362 430
rect 7478 400 8370 430
rect 8486 400 9378 430
rect 9494 400 10386 430
rect 10502 400 11394 430
rect 11510 400 12402 430
rect 12518 400 13410 430
rect 13526 400 14418 430
rect 14534 400 15426 430
rect 15542 400 16434 430
rect 16550 400 17442 430
rect 17558 400 18450 430
rect 18566 400 19458 430
rect 19574 400 20466 430
rect 20582 400 21474 430
rect 21590 400 22482 430
rect 22598 400 23490 430
rect 23606 400 24122 430
<< metal3 >>
rect 0 23744 400 23800
rect 24600 23184 25000 23240
rect 0 22960 400 23016
rect 0 22176 400 22232
rect 0 21392 400 21448
rect 0 20608 400 20664
rect 24600 20496 25000 20552
rect 0 19824 400 19880
rect 0 19040 400 19096
rect 0 18256 400 18312
rect 24600 17808 25000 17864
rect 0 17472 400 17528
rect 0 16688 400 16744
rect 0 15904 400 15960
rect 0 15120 400 15176
rect 24600 15120 25000 15176
rect 0 14336 400 14392
rect 0 13552 400 13608
rect 0 12768 400 12824
rect 24600 12432 25000 12488
rect 0 11984 400 12040
rect 0 11200 400 11256
rect 0 10416 400 10472
rect 24600 9744 25000 9800
rect 0 9632 400 9688
rect 0 8848 400 8904
rect 0 8064 400 8120
rect 0 7280 400 7336
rect 24600 7056 25000 7112
rect 0 6496 400 6552
rect 0 5712 400 5768
rect 0 4928 400 4984
rect 24600 4368 25000 4424
rect 0 4144 400 4200
rect 0 3360 400 3416
rect 0 2576 400 2632
rect 0 1792 400 1848
rect 24600 1680 25000 1736
rect 0 1008 400 1064
<< obsm3 >>
rect 430 23714 24600 23786
rect 400 23270 24600 23714
rect 400 23154 24570 23270
rect 400 23046 24600 23154
rect 430 22930 24600 23046
rect 400 22262 24600 22930
rect 430 22146 24600 22262
rect 400 21478 24600 22146
rect 430 21362 24600 21478
rect 400 20694 24600 21362
rect 430 20582 24600 20694
rect 430 20578 24570 20582
rect 400 20466 24570 20578
rect 400 19910 24600 20466
rect 430 19794 24600 19910
rect 400 19126 24600 19794
rect 430 19010 24600 19126
rect 400 18342 24600 19010
rect 430 18226 24600 18342
rect 400 17894 24600 18226
rect 400 17778 24570 17894
rect 400 17558 24600 17778
rect 430 17442 24600 17558
rect 400 16774 24600 17442
rect 430 16658 24600 16774
rect 400 15990 24600 16658
rect 430 15874 24600 15990
rect 400 15206 24600 15874
rect 430 15090 24570 15206
rect 400 14422 24600 15090
rect 430 14306 24600 14422
rect 400 13638 24600 14306
rect 430 13522 24600 13638
rect 400 12854 24600 13522
rect 430 12738 24600 12854
rect 400 12518 24600 12738
rect 400 12402 24570 12518
rect 400 12070 24600 12402
rect 430 11954 24600 12070
rect 400 11286 24600 11954
rect 430 11170 24600 11286
rect 400 10502 24600 11170
rect 430 10386 24600 10502
rect 400 9830 24600 10386
rect 400 9718 24570 9830
rect 430 9714 24570 9718
rect 430 9602 24600 9714
rect 400 8934 24600 9602
rect 430 8818 24600 8934
rect 400 8150 24600 8818
rect 430 8034 24600 8150
rect 400 7366 24600 8034
rect 430 7250 24600 7366
rect 400 7142 24600 7250
rect 400 7026 24570 7142
rect 400 6582 24600 7026
rect 430 6466 24600 6582
rect 400 5798 24600 6466
rect 430 5682 24600 5798
rect 400 5014 24600 5682
rect 430 4898 24600 5014
rect 400 4454 24600 4898
rect 400 4338 24570 4454
rect 400 4230 24600 4338
rect 430 4114 24600 4230
rect 400 3446 24600 4114
rect 430 3330 24600 3446
rect 400 2662 24600 3330
rect 430 2546 24600 2662
rect 400 1878 24600 2546
rect 430 1766 24600 1878
rect 430 1762 24570 1766
rect 400 1650 24570 1762
rect 400 1094 24600 1650
rect 430 1022 24600 1094
<< metal4 >>
rect 2224 1538 2384 23158
rect 9904 1538 10064 23158
rect 17584 1538 17744 23158
<< obsm4 >>
rect 2478 4769 9874 22559
rect 10094 4769 17234 22559
<< labels >>
rlabel metal3 s 24600 15120 25000 15176 6 DAC_clk
port 1 nsew signal input
rlabel metal3 s 24600 17808 25000 17864 6 DAC_d1
port 2 nsew signal input
rlabel metal3 s 24600 20496 25000 20552 6 DAC_d2
port 3 nsew signal input
rlabel metal3 s 24600 23184 25000 23240 6 DAC_le
port 4 nsew signal input
rlabel metal3 s 0 17472 400 17528 6 RXD
port 5 nsew signal output
rlabel metal3 s 0 16688 400 16744 6 TXD
port 6 nsew signal input
rlabel metal3 s 0 1008 400 1064 6 addr[0]
port 7 nsew signal input
rlabel metal3 s 0 1792 400 1848 6 addr[1]
port 8 nsew signal input
rlabel metal3 s 0 2576 400 2632 6 addr[2]
port 9 nsew signal input
rlabel metal3 s 0 3360 400 3416 6 addr[3]
port 10 nsew signal input
rlabel metal2 s 17472 0 17528 400 6 bus_cyc
port 11 nsew signal input
rlabel metal2 s 18480 0 18536 400 6 bus_we
port 12 nsew signal input
rlabel metal3 s 0 4144 400 4200 6 data_in[0]
port 13 nsew signal input
rlabel metal3 s 0 4928 400 4984 6 data_in[1]
port 14 nsew signal input
rlabel metal3 s 0 5712 400 5768 6 data_in[2]
port 15 nsew signal input
rlabel metal3 s 0 6496 400 6552 6 data_in[3]
port 16 nsew signal input
rlabel metal3 s 0 7280 400 7336 6 data_in[4]
port 17 nsew signal input
rlabel metal3 s 0 8064 400 8120 6 data_in[5]
port 18 nsew signal input
rlabel metal3 s 0 8848 400 8904 6 data_in[6]
port 19 nsew signal input
rlabel metal3 s 0 9632 400 9688 6 data_in[7]
port 20 nsew signal input
rlabel metal3 s 0 10416 400 10472 6 data_out[0]
port 21 nsew signal output
rlabel metal3 s 0 11200 400 11256 6 data_out[1]
port 22 nsew signal output
rlabel metal3 s 0 11984 400 12040 6 data_out[2]
port 23 nsew signal output
rlabel metal3 s 0 12768 400 12824 6 data_out[3]
port 24 nsew signal output
rlabel metal3 s 0 13552 400 13608 6 data_out[4]
port 25 nsew signal output
rlabel metal3 s 0 14336 400 14392 6 data_out[5]
port 26 nsew signal output
rlabel metal3 s 0 15120 400 15176 6 data_out[6]
port 27 nsew signal output
rlabel metal3 s 0 15904 400 15960 6 data_out[7]
port 28 nsew signal output
rlabel metal2 s 1344 24600 1400 25000 6 io_in[0]
port 29 nsew signal input
rlabel metal2 s 8064 24600 8120 25000 6 io_in[10]
port 30 nsew signal input
rlabel metal2 s 8736 24600 8792 25000 6 io_in[11]
port 31 nsew signal input
rlabel metal2 s 9408 24600 9464 25000 6 io_in[12]
port 32 nsew signal input
rlabel metal2 s 10080 24600 10136 25000 6 io_in[13]
port 33 nsew signal input
rlabel metal2 s 10752 24600 10808 25000 6 io_in[14]
port 34 nsew signal input
rlabel metal2 s 11424 24600 11480 25000 6 io_in[15]
port 35 nsew signal input
rlabel metal2 s 2016 24600 2072 25000 6 io_in[1]
port 36 nsew signal input
rlabel metal2 s 2688 24600 2744 25000 6 io_in[2]
port 37 nsew signal input
rlabel metal2 s 3360 24600 3416 25000 6 io_in[3]
port 38 nsew signal input
rlabel metal2 s 4032 24600 4088 25000 6 io_in[4]
port 39 nsew signal input
rlabel metal2 s 4704 24600 4760 25000 6 io_in[5]
port 40 nsew signal input
rlabel metal2 s 5376 24600 5432 25000 6 io_in[6]
port 41 nsew signal input
rlabel metal2 s 6048 24600 6104 25000 6 io_in[7]
port 42 nsew signal input
rlabel metal2 s 6720 24600 6776 25000 6 io_in[8]
port 43 nsew signal input
rlabel metal2 s 7392 24600 7448 25000 6 io_in[9]
port 44 nsew signal input
rlabel metal2 s 1344 0 1400 400 6 io_oeb[0]
port 45 nsew signal output
rlabel metal2 s 11424 0 11480 400 6 io_oeb[10]
port 46 nsew signal output
rlabel metal2 s 12432 0 12488 400 6 io_oeb[11]
port 47 nsew signal output
rlabel metal2 s 13440 0 13496 400 6 io_oeb[12]
port 48 nsew signal output
rlabel metal2 s 14448 0 14504 400 6 io_oeb[13]
port 49 nsew signal output
rlabel metal2 s 15456 0 15512 400 6 io_oeb[14]
port 50 nsew signal output
rlabel metal2 s 16464 0 16520 400 6 io_oeb[15]
port 51 nsew signal output
rlabel metal2 s 2352 0 2408 400 6 io_oeb[1]
port 52 nsew signal output
rlabel metal2 s 3360 0 3416 400 6 io_oeb[2]
port 53 nsew signal output
rlabel metal2 s 4368 0 4424 400 6 io_oeb[3]
port 54 nsew signal output
rlabel metal2 s 5376 0 5432 400 6 io_oeb[4]
port 55 nsew signal output
rlabel metal2 s 6384 0 6440 400 6 io_oeb[5]
port 56 nsew signal output
rlabel metal2 s 7392 0 7448 400 6 io_oeb[6]
port 57 nsew signal output
rlabel metal2 s 8400 0 8456 400 6 io_oeb[7]
port 58 nsew signal output
rlabel metal2 s 9408 0 9464 400 6 io_oeb[8]
port 59 nsew signal output
rlabel metal2 s 10416 0 10472 400 6 io_oeb[9]
port 60 nsew signal output
rlabel metal2 s 12096 24600 12152 25000 6 io_out[0]
port 61 nsew signal output
rlabel metal2 s 18816 24600 18872 25000 6 io_out[10]
port 62 nsew signal output
rlabel metal2 s 19488 24600 19544 25000 6 io_out[11]
port 63 nsew signal output
rlabel metal2 s 20160 24600 20216 25000 6 io_out[12]
port 64 nsew signal output
rlabel metal2 s 20832 24600 20888 25000 6 io_out[13]
port 65 nsew signal output
rlabel metal2 s 21504 24600 21560 25000 6 io_out[14]
port 66 nsew signal output
rlabel metal2 s 22176 24600 22232 25000 6 io_out[15]
port 67 nsew signal output
rlabel metal2 s 12768 24600 12824 25000 6 io_out[1]
port 68 nsew signal output
rlabel metal2 s 13440 24600 13496 25000 6 io_out[2]
port 69 nsew signal output
rlabel metal2 s 14112 24600 14168 25000 6 io_out[3]
port 70 nsew signal output
rlabel metal2 s 14784 24600 14840 25000 6 io_out[4]
port 71 nsew signal output
rlabel metal2 s 15456 24600 15512 25000 6 io_out[5]
port 72 nsew signal output
rlabel metal2 s 16128 24600 16184 25000 6 io_out[6]
port 73 nsew signal output
rlabel metal2 s 16800 24600 16856 25000 6 io_out[7]
port 74 nsew signal output
rlabel metal2 s 17472 24600 17528 25000 6 io_out[8]
port 75 nsew signal output
rlabel metal2 s 18144 24600 18200 25000 6 io_out[9]
port 76 nsew signal output
rlabel metal2 s 19488 0 19544 400 6 irq0
port 77 nsew signal output
rlabel metal2 s 20496 0 20552 400 6 irq6
port 78 nsew signal output
rlabel metal2 s 21504 0 21560 400 6 irq7
port 79 nsew signal output
rlabel metal3 s 0 18256 400 18312 6 la_data_out[0]
port 80 nsew signal output
rlabel metal3 s 0 19040 400 19096 6 la_data_out[1]
port 81 nsew signal output
rlabel metal3 s 0 19824 400 19880 6 la_data_out[2]
port 82 nsew signal output
rlabel metal3 s 0 20608 400 20664 6 la_data_out[3]
port 83 nsew signal output
rlabel metal3 s 0 21392 400 21448 6 la_data_out[4]
port 84 nsew signal output
rlabel metal3 s 0 22176 400 22232 6 la_data_out[5]
port 85 nsew signal output
rlabel metal3 s 0 22960 400 23016 6 la_data_out[6]
port 86 nsew signal output
rlabel metal3 s 0 23744 400 23800 6 la_data_out[7]
port 87 nsew signal output
rlabel metal3 s 24600 7056 25000 7112 6 pwm0
port 88 nsew signal input
rlabel metal3 s 24600 9744 25000 9800 6 pwm1
port 89 nsew signal input
rlabel metal3 s 24600 12432 25000 12488 6 pwm2
port 90 nsew signal input
rlabel metal2 s 23520 0 23576 400 6 rst
port 91 nsew signal input
rlabel metal2 s 22848 24600 22904 25000 6 tmr0_clk
port 92 nsew signal output
rlabel metal3 s 24600 1680 25000 1736 6 tmr0_o
port 93 nsew signal input
rlabel metal2 s 23520 24600 23576 25000 6 tmr1_clk
port 94 nsew signal output
rlabel metal3 s 24600 4368 25000 4424 6 tmr1_o
port 95 nsew signal input
rlabel metal4 s 2224 1538 2384 23158 6 vdd
port 96 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 23158 6 vdd
port 96 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 23158 6 vss
port 97 nsew ground bidirectional
rlabel metal2 s 22512 0 22568 400 6 wb_clk_i
port 98 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 25000 25000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 1426344
string GDS_FILE /run/media/tholin/fbc90f8f-67e9-406d-9872-54f02ad6a2d8/AS2650/openlane/gpios/runs/23_11_20_21_39/results/signoff/gpios.magic.gds
string GDS_START 217822
<< end >>

